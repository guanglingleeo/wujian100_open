/*
Copyright (c) 2019 Alibaba Group Holding Limited

Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation files (the "Software"), to deal in the Software without restriction, including without limitation the rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the Software is furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.

*/
module ahb_matrix_7_12_arb(
  hclk,
  hresetn,
  m0_latch_cmd,
  m0_nor_hready,
  m0_s0_cmd_cur,
  m0_s0_cmd_last,
  m0_s0_data,
  m0_s0_req,
  m0_s10_cmd_cur,
  m0_s10_cmd_last,
  m0_s10_data,
  m0_s10_req,
  m0_s11_cmd_cur,
  m0_s11_cmd_last,
  m0_s11_data,
  m0_s11_req,
  m0_s1_cmd_cur,
  m0_s1_cmd_last,
  m0_s1_data,
  m0_s1_req,
  m0_s2_cmd_cur,
  m0_s2_cmd_last,
  m0_s2_data,
  m0_s2_req,
  m0_s3_cmd_cur,
  m0_s3_cmd_last,
  m0_s3_data,
  m0_s3_req,
  m0_s4_cmd_cur,
  m0_s4_cmd_last,
  m0_s4_data,
  m0_s4_req,
  m0_s5_cmd_cur,
  m0_s5_cmd_last,
  m0_s5_data,
  m0_s5_req,
  m0_s6_cmd_cur,
  m0_s6_cmd_last,
  m0_s6_data,
  m0_s6_req,
  m0_s7_cmd_cur,
  m0_s7_cmd_last,
  m0_s7_data,
  m0_s7_req,
  m0_s8_cmd_cur,
  m0_s8_cmd_last,
  m0_s8_data,
  m0_s8_req,
  m0_s9_cmd_cur,
  m0_s9_cmd_last,
  m0_s9_data,
  m0_s9_req,
  m1_latch_cmd,
  m1_nor_hready,
  m1_s0_cmd_cur,
  m1_s0_cmd_last,
  m1_s0_data,
  m1_s0_req,
  m1_s10_cmd_cur,
  m1_s10_cmd_last,
  m1_s10_data,
  m1_s10_req,
  m1_s11_cmd_cur,
  m1_s11_cmd_last,
  m1_s11_data,
  m1_s11_req,
  m1_s1_cmd_cur,
  m1_s1_cmd_last,
  m1_s1_data,
  m1_s1_req,
  m1_s2_cmd_cur,
  m1_s2_cmd_last,
  m1_s2_data,
  m1_s2_req,
  m1_s3_cmd_cur,
  m1_s3_cmd_last,
  m1_s3_data,
  m1_s3_req,
  m1_s4_cmd_cur,
  m1_s4_cmd_last,
  m1_s4_data,
  m1_s4_req,
  m1_s5_cmd_cur,
  m1_s5_cmd_last,
  m1_s5_data,
  m1_s5_req,
  m1_s6_cmd_cur,
  m1_s6_cmd_last,
  m1_s6_data,
  m1_s6_req,
  m1_s7_cmd_cur,
  m1_s7_cmd_last,
  m1_s7_data,
  m1_s7_req,
  m1_s8_cmd_cur,
  m1_s8_cmd_last,
  m1_s8_data,
  m1_s8_req,
  m1_s9_cmd_cur,
  m1_s9_cmd_last,
  m1_s9_data,
  m1_s9_req,
  m2_latch_cmd,
  m2_nor_hready,
  m2_s0_cmd_cur,
  m2_s0_cmd_last,
  m2_s0_data,
  m2_s0_req,
  m2_s10_cmd_cur,
  m2_s10_cmd_last,
  m2_s10_data,
  m2_s10_req,
  m2_s11_cmd_cur,
  m2_s11_cmd_last,
  m2_s11_data,
  m2_s11_req,
  m2_s1_cmd_cur,
  m2_s1_cmd_last,
  m2_s1_data,
  m2_s1_req,
  m2_s2_cmd_cur,
  m2_s2_cmd_last,
  m2_s2_data,
  m2_s2_req,
  m2_s3_cmd_cur,
  m2_s3_cmd_last,
  m2_s3_data,
  m2_s3_req,
  m2_s4_cmd_cur,
  m2_s4_cmd_last,
  m2_s4_data,
  m2_s4_req,
  m2_s5_cmd_cur,
  m2_s5_cmd_last,
  m2_s5_data,
  m2_s5_req,
  m2_s6_cmd_cur,
  m2_s6_cmd_last,
  m2_s6_data,
  m2_s6_req,
  m2_s7_cmd_cur,
  m2_s7_cmd_last,
  m2_s7_data,
  m2_s7_req,
  m2_s8_cmd_cur,
  m2_s8_cmd_last,
  m2_s8_data,
  m2_s8_req,
  m2_s9_cmd_cur,
  m2_s9_cmd_last,
  m2_s9_data,
  m2_s9_req,
  m3_latch_cmd,
  m3_nor_hready,
  m3_s0_cmd_cur,
  m3_s0_cmd_last,
  m3_s0_data,
  m3_s0_req,
  m3_s10_cmd_cur,
  m3_s10_cmd_last,
  m3_s10_data,
  m3_s10_req,
  m3_s11_cmd_cur,
  m3_s11_cmd_last,
  m3_s11_data,
  m3_s11_req,
  m3_s1_cmd_cur,
  m3_s1_cmd_last,
  m3_s1_data,
  m3_s1_req,
  m3_s2_cmd_cur,
  m3_s2_cmd_last,
  m3_s2_data,
  m3_s2_req,
  m3_s3_cmd_cur,
  m3_s3_cmd_last,
  m3_s3_data,
  m3_s3_req,
  m3_s4_cmd_cur,
  m3_s4_cmd_last,
  m3_s4_data,
  m3_s4_req,
  m3_s5_cmd_cur,
  m3_s5_cmd_last,
  m3_s5_data,
  m3_s5_req,
  m3_s6_cmd_cur,
  m3_s6_cmd_last,
  m3_s6_data,
  m3_s6_req,
  m3_s7_cmd_cur,
  m3_s7_cmd_last,
  m3_s7_data,
  m3_s7_req,
  m3_s8_cmd_cur,
  m3_s8_cmd_last,
  m3_s8_data,
  m3_s8_req,
  m3_s9_cmd_cur,
  m3_s9_cmd_last,
  m3_s9_data,
  m3_s9_req,
  m4_latch_cmd,
  m4_nor_hready,
  m4_s0_cmd_cur,
  m4_s0_cmd_last,
  m4_s0_data,
  m4_s0_req,
  m4_s10_cmd_cur,
  m4_s10_cmd_last,
  m4_s10_data,
  m4_s10_req,
  m4_s11_cmd_cur,
  m4_s11_cmd_last,
  m4_s11_data,
  m4_s11_req,
  m4_s1_cmd_cur,
  m4_s1_cmd_last,
  m4_s1_data,
  m4_s1_req,
  m4_s2_cmd_cur,
  m4_s2_cmd_last,
  m4_s2_data,
  m4_s2_req,
  m4_s3_cmd_cur,
  m4_s3_cmd_last,
  m4_s3_data,
  m4_s3_req,
  m4_s4_cmd_cur,
  m4_s4_cmd_last,
  m4_s4_data,
  m4_s4_req,
  m4_s5_cmd_cur,
  m4_s5_cmd_last,
  m4_s5_data,
  m4_s5_req,
  m4_s6_cmd_cur,
  m4_s6_cmd_last,
  m4_s6_data,
  m4_s6_req,
  m4_s7_cmd_cur,
  m4_s7_cmd_last,
  m4_s7_data,
  m4_s7_req,
  m4_s8_cmd_cur,
  m4_s8_cmd_last,
  m4_s8_data,
  m4_s8_req,
  m4_s9_cmd_cur,
  m4_s9_cmd_last,
  m4_s9_data,
  m4_s9_req,
  m5_latch_cmd,
  m5_nor_hready,
  m5_s0_cmd_cur,
  m5_s0_cmd_last,
  m5_s0_data,
  m5_s0_req,
  m5_s10_cmd_cur,
  m5_s10_cmd_last,
  m5_s10_data,
  m5_s10_req,
  m5_s11_cmd_cur,
  m5_s11_cmd_last,
  m5_s11_data,
  m5_s11_req,
  m5_s1_cmd_cur,
  m5_s1_cmd_last,
  m5_s1_data,
  m5_s1_req,
  m5_s2_cmd_cur,
  m5_s2_cmd_last,
  m5_s2_data,
  m5_s2_req,
  m5_s3_cmd_cur,
  m5_s3_cmd_last,
  m5_s3_data,
  m5_s3_req,
  m5_s4_cmd_cur,
  m5_s4_cmd_last,
  m5_s4_data,
  m5_s4_req,
  m5_s5_cmd_cur,
  m5_s5_cmd_last,
  m5_s5_data,
  m5_s5_req,
  m5_s6_cmd_cur,
  m5_s6_cmd_last,
  m5_s6_data,
  m5_s6_req,
  m5_s7_cmd_cur,
  m5_s7_cmd_last,
  m5_s7_data,
  m5_s7_req,
  m5_s8_cmd_cur,
  m5_s8_cmd_last,
  m5_s8_data,
  m5_s8_req,
  m5_s9_cmd_cur,
  m5_s9_cmd_last,
  m5_s9_data,
  m5_s9_req,
  m6_latch_cmd,
  m6_nor_hready,
  m6_s0_cmd_cur,
  m6_s0_cmd_last,
  m6_s0_data,
  m6_s0_req,
  m6_s10_cmd_cur,
  m6_s10_cmd_last,
  m6_s10_data,
  m6_s10_req,
  m6_s11_cmd_cur,
  m6_s11_cmd_last,
  m6_s11_data,
  m6_s11_req,
  m6_s1_cmd_cur,
  m6_s1_cmd_last,
  m6_s1_data,
  m6_s1_req,
  m6_s2_cmd_cur,
  m6_s2_cmd_last,
  m6_s2_data,
  m6_s2_req,
  m6_s3_cmd_cur,
  m6_s3_cmd_last,
  m6_s3_data,
  m6_s3_req,
  m6_s4_cmd_cur,
  m6_s4_cmd_last,
  m6_s4_data,
  m6_s4_req,
  m6_s5_cmd_cur,
  m6_s5_cmd_last,
  m6_s5_data,
  m6_s5_req,
  m6_s6_cmd_cur,
  m6_s6_cmd_last,
  m6_s6_data,
  m6_s6_req,
  m6_s7_cmd_cur,
  m6_s7_cmd_last,
  m6_s7_data,
  m6_s7_req,
  m6_s8_cmd_cur,
  m6_s8_cmd_last,
  m6_s8_data,
  m6_s8_req,
  m6_s9_cmd_cur,
  m6_s9_cmd_last,
  m6_s9_data,
  m6_s9_req,
  s0_hready,
  s0_req,
  s10_hready,
  s10_req,
  s11_hready,
  s11_req,
  s1_hready,
  s1_req,
  s2_hready,
  s2_req,
  s3_hready,
  s3_req,
  s4_hready,
  s4_req,
  s5_hready,
  s5_req,
  s6_hready,
  s6_req,
  s7_hready,
  s7_req,
  s8_hready,
  s8_req,
  s9_hready,
  s9_req
);
input           hclk;               
input           hresetn;            
input           m0_s0_req;          
input           m0_s10_req;         
input           m0_s11_req;         
input           m0_s1_req;          
input           m0_s2_req;          
input           m0_s3_req;          
input           m0_s4_req;          
input           m0_s5_req;          
input           m0_s6_req;          
input           m0_s7_req;          
input           m0_s8_req;          
input           m0_s9_req;          
input           m1_s0_req;          
input           m1_s10_req;         
input           m1_s11_req;         
input           m1_s1_req;          
input           m1_s2_req;          
input           m1_s3_req;          
input           m1_s4_req;          
input           m1_s5_req;          
input           m1_s6_req;          
input           m1_s7_req;          
input           m1_s8_req;          
input           m1_s9_req;          
input           m2_s0_req;          
input           m2_s10_req;         
input           m2_s11_req;         
input           m2_s1_req;          
input           m2_s2_req;          
input           m2_s3_req;          
input           m2_s4_req;          
input           m2_s5_req;          
input           m2_s6_req;          
input           m2_s7_req;          
input           m2_s8_req;          
input           m2_s9_req;          
input           m3_s0_req;          
input           m3_s10_req;         
input           m3_s11_req;         
input           m3_s1_req;          
input           m3_s2_req;          
input           m3_s3_req;          
input           m3_s4_req;          
input           m3_s5_req;          
input           m3_s6_req;          
input           m3_s7_req;          
input           m3_s8_req;          
input           m3_s9_req;          
input           m4_s0_req;          
input           m4_s10_req;         
input           m4_s11_req;         
input           m4_s1_req;          
input           m4_s2_req;          
input           m4_s3_req;          
input           m4_s4_req;          
input           m4_s5_req;          
input           m4_s6_req;          
input           m4_s7_req;          
input           m4_s8_req;          
input           m4_s9_req;          
input           m5_s0_req;          
input           m5_s10_req;         
input           m5_s11_req;         
input           m5_s1_req;          
input           m5_s2_req;          
input           m5_s3_req;          
input           m5_s4_req;          
input           m5_s5_req;          
input           m5_s6_req;          
input           m5_s7_req;          
input           m5_s8_req;          
input           m5_s9_req;          
input           m6_s0_req;          
input           m6_s10_req;         
input           m6_s11_req;         
input           m6_s1_req;          
input           m6_s2_req;          
input           m6_s3_req;          
input           m6_s4_req;          
input           m6_s5_req;          
input           m6_s6_req;          
input           m6_s7_req;          
input           m6_s8_req;          
input           m6_s9_req;          
input           s0_hready;          
input   [6 :0]  s0_req;             
input           s10_hready;         
input   [6 :0]  s10_req;            
input           s11_hready;         
input   [6 :0]  s11_req;            
input           s1_hready;          
input   [6 :0]  s1_req;             
input           s2_hready;          
input   [6 :0]  s2_req;             
input           s3_hready;          
input   [6 :0]  s3_req;             
input           s4_hready;          
input   [6 :0]  s4_req;             
input           s5_hready;          
input   [6 :0]  s5_req;             
input           s6_hready;          
input   [6 :0]  s6_req;             
input           s7_hready;          
input   [6 :0]  s7_req;             
input           s8_hready;          
input   [6 :0]  s8_req;             
input           s9_hready;          
input   [6 :0]  s9_req;             
output          m0_latch_cmd;       
output          m0_nor_hready;      
output          m0_s0_cmd_cur;      
output          m0_s0_cmd_last;     
output          m0_s0_data;         
output          m0_s10_cmd_cur;     
output          m0_s10_cmd_last;    
output          m0_s10_data;        
output          m0_s11_cmd_cur;     
output          m0_s11_cmd_last;    
output          m0_s11_data;        
output          m0_s1_cmd_cur;      
output          m0_s1_cmd_last;     
output          m0_s1_data;         
output          m0_s2_cmd_cur;      
output          m0_s2_cmd_last;     
output          m0_s2_data;         
output          m0_s3_cmd_cur;      
output          m0_s3_cmd_last;     
output          m0_s3_data;         
output          m0_s4_cmd_cur;      
output          m0_s4_cmd_last;     
output          m0_s4_data;         
output          m0_s5_cmd_cur;      
output          m0_s5_cmd_last;     
output          m0_s5_data;         
output          m0_s6_cmd_cur;      
output          m0_s6_cmd_last;     
output          m0_s6_data;         
output          m0_s7_cmd_cur;      
output          m0_s7_cmd_last;     
output          m0_s7_data;         
output          m0_s8_cmd_cur;      
output          m0_s8_cmd_last;     
output          m0_s8_data;         
output          m0_s9_cmd_cur;      
output          m0_s9_cmd_last;     
output          m0_s9_data;         
output          m1_latch_cmd;       
output          m1_nor_hready;      
output          m1_s0_cmd_cur;      
output          m1_s0_cmd_last;     
output          m1_s0_data;         
output          m1_s10_cmd_cur;     
output          m1_s10_cmd_last;    
output          m1_s10_data;        
output          m1_s11_cmd_cur;     
output          m1_s11_cmd_last;    
output          m1_s11_data;        
output          m1_s1_cmd_cur;      
output          m1_s1_cmd_last;     
output          m1_s1_data;         
output          m1_s2_cmd_cur;      
output          m1_s2_cmd_last;     
output          m1_s2_data;         
output          m1_s3_cmd_cur;      
output          m1_s3_cmd_last;     
output          m1_s3_data;         
output          m1_s4_cmd_cur;      
output          m1_s4_cmd_last;     
output          m1_s4_data;         
output          m1_s5_cmd_cur;      
output          m1_s5_cmd_last;     
output          m1_s5_data;         
output          m1_s6_cmd_cur;      
output          m1_s6_cmd_last;     
output          m1_s6_data;         
output          m1_s7_cmd_cur;      
output          m1_s7_cmd_last;     
output          m1_s7_data;         
output          m1_s8_cmd_cur;      
output          m1_s8_cmd_last;     
output          m1_s8_data;         
output          m1_s9_cmd_cur;      
output          m1_s9_cmd_last;     
output          m1_s9_data;         
output          m2_latch_cmd;       
output          m2_nor_hready;      
output          m2_s0_cmd_cur;      
output          m2_s0_cmd_last;     
output          m2_s0_data;         
output          m2_s10_cmd_cur;     
output          m2_s10_cmd_last;    
output          m2_s10_data;        
output          m2_s11_cmd_cur;     
output          m2_s11_cmd_last;    
output          m2_s11_data;        
output          m2_s1_cmd_cur;      
output          m2_s1_cmd_last;     
output          m2_s1_data;         
output          m2_s2_cmd_cur;      
output          m2_s2_cmd_last;     
output          m2_s2_data;         
output          m2_s3_cmd_cur;      
output          m2_s3_cmd_last;     
output          m2_s3_data;         
output          m2_s4_cmd_cur;      
output          m2_s4_cmd_last;     
output          m2_s4_data;         
output          m2_s5_cmd_cur;      
output          m2_s5_cmd_last;     
output          m2_s5_data;         
output          m2_s6_cmd_cur;      
output          m2_s6_cmd_last;     
output          m2_s6_data;         
output          m2_s7_cmd_cur;      
output          m2_s7_cmd_last;     
output          m2_s7_data;         
output          m2_s8_cmd_cur;      
output          m2_s8_cmd_last;     
output          m2_s8_data;         
output          m2_s9_cmd_cur;      
output          m2_s9_cmd_last;     
output          m2_s9_data;         
output          m3_latch_cmd;       
output          m3_nor_hready;      
output          m3_s0_cmd_cur;      
output          m3_s0_cmd_last;     
output          m3_s0_data;         
output          m3_s10_cmd_cur;     
output          m3_s10_cmd_last;    
output          m3_s10_data;        
output          m3_s11_cmd_cur;     
output          m3_s11_cmd_last;    
output          m3_s11_data;        
output          m3_s1_cmd_cur;      
output          m3_s1_cmd_last;     
output          m3_s1_data;         
output          m3_s2_cmd_cur;      
output          m3_s2_cmd_last;     
output          m3_s2_data;         
output          m3_s3_cmd_cur;      
output          m3_s3_cmd_last;     
output          m3_s3_data;         
output          m3_s4_cmd_cur;      
output          m3_s4_cmd_last;     
output          m3_s4_data;         
output          m3_s5_cmd_cur;      
output          m3_s5_cmd_last;     
output          m3_s5_data;         
output          m3_s6_cmd_cur;      
output          m3_s6_cmd_last;     
output          m3_s6_data;         
output          m3_s7_cmd_cur;      
output          m3_s7_cmd_last;     
output          m3_s7_data;         
output          m3_s8_cmd_cur;      
output          m3_s8_cmd_last;     
output          m3_s8_data;         
output          m3_s9_cmd_cur;      
output          m3_s9_cmd_last;     
output          m3_s9_data;         
output          m4_latch_cmd;       
output          m4_nor_hready;      
output          m4_s0_cmd_cur;      
output          m4_s0_cmd_last;     
output          m4_s0_data;         
output          m4_s10_cmd_cur;     
output          m4_s10_cmd_last;    
output          m4_s10_data;        
output          m4_s11_cmd_cur;     
output          m4_s11_cmd_last;    
output          m4_s11_data;        
output          m4_s1_cmd_cur;      
output          m4_s1_cmd_last;     
output          m4_s1_data;         
output          m4_s2_cmd_cur;      
output          m4_s2_cmd_last;     
output          m4_s2_data;         
output          m4_s3_cmd_cur;      
output          m4_s3_cmd_last;     
output          m4_s3_data;         
output          m4_s4_cmd_cur;      
output          m4_s4_cmd_last;     
output          m4_s4_data;         
output          m4_s5_cmd_cur;      
output          m4_s5_cmd_last;     
output          m4_s5_data;         
output          m4_s6_cmd_cur;      
output          m4_s6_cmd_last;     
output          m4_s6_data;         
output          m4_s7_cmd_cur;      
output          m4_s7_cmd_last;     
output          m4_s7_data;         
output          m4_s8_cmd_cur;      
output          m4_s8_cmd_last;     
output          m4_s8_data;         
output          m4_s9_cmd_cur;      
output          m4_s9_cmd_last;     
output          m4_s9_data;         
output          m5_latch_cmd;       
output          m5_nor_hready;      
output          m5_s0_cmd_cur;      
output          m5_s0_cmd_last;     
output          m5_s0_data;         
output          m5_s10_cmd_cur;     
output          m5_s10_cmd_last;    
output          m5_s10_data;        
output          m5_s11_cmd_cur;     
output          m5_s11_cmd_last;    
output          m5_s11_data;        
output          m5_s1_cmd_cur;      
output          m5_s1_cmd_last;     
output          m5_s1_data;         
output          m5_s2_cmd_cur;      
output          m5_s2_cmd_last;     
output          m5_s2_data;         
output          m5_s3_cmd_cur;      
output          m5_s3_cmd_last;     
output          m5_s3_data;         
output          m5_s4_cmd_cur;      
output          m5_s4_cmd_last;     
output          m5_s4_data;         
output          m5_s5_cmd_cur;      
output          m5_s5_cmd_last;     
output          m5_s5_data;         
output          m5_s6_cmd_cur;      
output          m5_s6_cmd_last;     
output          m5_s6_data;         
output          m5_s7_cmd_cur;      
output          m5_s7_cmd_last;     
output          m5_s7_data;         
output          m5_s8_cmd_cur;      
output          m5_s8_cmd_last;     
output          m5_s8_data;         
output          m5_s9_cmd_cur;      
output          m5_s9_cmd_last;     
output          m5_s9_data;         
output          m6_latch_cmd;       
output          m6_nor_hready;      
output          m6_s0_cmd_cur;      
output          m6_s0_cmd_last;     
output          m6_s0_data;         
output          m6_s10_cmd_cur;     
output          m6_s10_cmd_last;    
output          m6_s10_data;        
output          m6_s11_cmd_cur;     
output          m6_s11_cmd_last;    
output          m6_s11_data;        
output          m6_s1_cmd_cur;      
output          m6_s1_cmd_last;     
output          m6_s1_data;         
output          m6_s2_cmd_cur;      
output          m6_s2_cmd_last;     
output          m6_s2_data;         
output          m6_s3_cmd_cur;      
output          m6_s3_cmd_last;     
output          m6_s3_data;         
output          m6_s4_cmd_cur;      
output          m6_s4_cmd_last;     
output          m6_s4_data;         
output          m6_s5_cmd_cur;      
output          m6_s5_cmd_last;     
output          m6_s5_data;         
output          m6_s6_cmd_cur;      
output          m6_s6_cmd_last;     
output          m6_s6_data;         
output          m6_s7_cmd_cur;      
output          m6_s7_cmd_last;     
output          m6_s7_data;         
output          m6_s8_cmd_cur;      
output          m6_s8_cmd_last;     
output          m6_s8_data;         
output          m6_s9_cmd_cur;      
output          m6_s9_cmd_last;     
output          m6_s9_data;         
reg     [48:0]  m0_cur_st;          
reg             m0_latch_cmd;       
reg             m0_nor_hready;      
reg     [48:0]  m0_nxt_st;          
reg             m0_s0_cmd_cur;      
reg             m0_s0_cmd_last;     
reg             m0_s0_data;         
reg             m0_s0_req_pend_tmp; 
reg             m0_s10_cmd_cur;     
reg             m0_s10_cmd_last;    
reg             m0_s10_data;        
reg             m0_s10_req_pend_tmp; 
reg             m0_s11_cmd_cur;     
reg             m0_s11_cmd_last;    
reg             m0_s11_data;        
reg             m0_s11_req_pend_tmp; 
reg             m0_s1_cmd_cur;      
reg             m0_s1_cmd_last;     
reg             m0_s1_data;         
reg             m0_s1_req_pend_tmp; 
reg             m0_s2_cmd_cur;      
reg             m0_s2_cmd_last;     
reg             m0_s2_data;         
reg             m0_s2_req_pend_tmp; 
reg             m0_s3_cmd_cur;      
reg             m0_s3_cmd_last;     
reg             m0_s3_data;         
reg             m0_s3_req_pend_tmp; 
reg             m0_s4_cmd_cur;      
reg             m0_s4_cmd_last;     
reg             m0_s4_data;         
reg             m0_s4_req_pend_tmp; 
reg             m0_s5_cmd_cur;      
reg             m0_s5_cmd_last;     
reg             m0_s5_data;         
reg             m0_s5_req_pend_tmp; 
reg             m0_s6_cmd_cur;      
reg             m0_s6_cmd_last;     
reg             m0_s6_data;         
reg             m0_s6_req_pend_tmp; 
reg             m0_s7_cmd_cur;      
reg             m0_s7_cmd_last;     
reg             m0_s7_data;         
reg             m0_s7_req_pend_tmp; 
reg             m0_s8_cmd_cur;      
reg             m0_s8_cmd_last;     
reg             m0_s8_data;         
reg             m0_s8_req_pend_tmp; 
reg             m0_s9_cmd_cur;      
reg             m0_s9_cmd_last;     
reg             m0_s9_data;         
reg             m0_s9_req_pend_tmp; 
reg     [48:0]  m1_cur_st;          
reg             m1_latch_cmd;       
reg             m1_nor_hready;      
reg     [48:0]  m1_nxt_st;          
reg             m1_s0_cmd_cur;      
reg             m1_s0_cmd_last;     
reg             m1_s0_data;         
reg             m1_s0_req_pend_tmp; 
reg             m1_s10_cmd_cur;     
reg             m1_s10_cmd_last;    
reg             m1_s10_data;        
reg             m1_s10_req_pend_tmp; 
reg             m1_s11_cmd_cur;     
reg             m1_s11_cmd_last;    
reg             m1_s11_data;        
reg             m1_s11_req_pend_tmp; 
reg             m1_s1_cmd_cur;      
reg             m1_s1_cmd_last;     
reg             m1_s1_data;         
reg             m1_s1_req_pend_tmp; 
reg             m1_s2_cmd_cur;      
reg             m1_s2_cmd_last;     
reg             m1_s2_data;         
reg             m1_s2_req_pend_tmp; 
reg             m1_s3_cmd_cur;      
reg             m1_s3_cmd_last;     
reg             m1_s3_data;         
reg             m1_s3_req_pend_tmp; 
reg             m1_s4_cmd_cur;      
reg             m1_s4_cmd_last;     
reg             m1_s4_data;         
reg             m1_s4_req_pend_tmp; 
reg             m1_s5_cmd_cur;      
reg             m1_s5_cmd_last;     
reg             m1_s5_data;         
reg             m1_s5_req_pend_tmp; 
reg             m1_s6_cmd_cur;      
reg             m1_s6_cmd_last;     
reg             m1_s6_data;         
reg             m1_s6_req_pend_tmp; 
reg             m1_s7_cmd_cur;      
reg             m1_s7_cmd_last;     
reg             m1_s7_data;         
reg             m1_s7_req_pend_tmp; 
reg             m1_s8_cmd_cur;      
reg             m1_s8_cmd_last;     
reg             m1_s8_data;         
reg             m1_s8_req_pend_tmp; 
reg             m1_s9_cmd_cur;      
reg             m1_s9_cmd_last;     
reg             m1_s9_data;         
reg             m1_s9_req_pend_tmp; 
reg     [48:0]  m2_cur_st;          
reg             m2_latch_cmd;       
reg             m2_nor_hready;      
reg     [48:0]  m2_nxt_st;          
reg             m2_s0_cmd_cur;      
reg             m2_s0_cmd_last;     
reg             m2_s0_data;         
reg             m2_s0_req_pend_tmp; 
reg             m2_s10_cmd_cur;     
reg             m2_s10_cmd_last;    
reg             m2_s10_data;        
reg             m2_s10_req_pend_tmp; 
reg             m2_s11_cmd_cur;     
reg             m2_s11_cmd_last;    
reg             m2_s11_data;        
reg             m2_s11_req_pend_tmp; 
reg             m2_s1_cmd_cur;      
reg             m2_s1_cmd_last;     
reg             m2_s1_data;         
reg             m2_s1_req_pend_tmp; 
reg             m2_s2_cmd_cur;      
reg             m2_s2_cmd_last;     
reg             m2_s2_data;         
reg             m2_s2_req_pend_tmp; 
reg             m2_s3_cmd_cur;      
reg             m2_s3_cmd_last;     
reg             m2_s3_data;         
reg             m2_s3_req_pend_tmp; 
reg             m2_s4_cmd_cur;      
reg             m2_s4_cmd_last;     
reg             m2_s4_data;         
reg             m2_s4_req_pend_tmp; 
reg             m2_s5_cmd_cur;      
reg             m2_s5_cmd_last;     
reg             m2_s5_data;         
reg             m2_s5_req_pend_tmp; 
reg             m2_s6_cmd_cur;      
reg             m2_s6_cmd_last;     
reg             m2_s6_data;         
reg             m2_s6_req_pend_tmp; 
reg             m2_s7_cmd_cur;      
reg             m2_s7_cmd_last;     
reg             m2_s7_data;         
reg             m2_s7_req_pend_tmp; 
reg             m2_s8_cmd_cur;      
reg             m2_s8_cmd_last;     
reg             m2_s8_data;         
reg             m2_s8_req_pend_tmp; 
reg             m2_s9_cmd_cur;      
reg             m2_s9_cmd_last;     
reg             m2_s9_data;         
reg             m2_s9_req_pend_tmp; 
reg     [48:0]  m3_cur_st;          
reg             m3_latch_cmd;       
reg             m3_nor_hready;      
reg     [48:0]  m3_nxt_st;          
reg             m3_s0_cmd_cur;      
reg             m3_s0_cmd_last;     
reg             m3_s0_data;         
reg             m3_s0_req_pend_tmp; 
reg             m3_s10_cmd_cur;     
reg             m3_s10_cmd_last;    
reg             m3_s10_data;        
reg             m3_s10_req_pend_tmp; 
reg             m3_s11_cmd_cur;     
reg             m3_s11_cmd_last;    
reg             m3_s11_data;        
reg             m3_s11_req_pend_tmp; 
reg             m3_s1_cmd_cur;      
reg             m3_s1_cmd_last;     
reg             m3_s1_data;         
reg             m3_s1_req_pend_tmp; 
reg             m3_s2_cmd_cur;      
reg             m3_s2_cmd_last;     
reg             m3_s2_data;         
reg             m3_s2_req_pend_tmp; 
reg             m3_s3_cmd_cur;      
reg             m3_s3_cmd_last;     
reg             m3_s3_data;         
reg             m3_s3_req_pend_tmp; 
reg             m3_s4_cmd_cur;      
reg             m3_s4_cmd_last;     
reg             m3_s4_data;         
reg             m3_s4_req_pend_tmp; 
reg             m3_s5_cmd_cur;      
reg             m3_s5_cmd_last;     
reg             m3_s5_data;         
reg             m3_s5_req_pend_tmp; 
reg             m3_s6_cmd_cur;      
reg             m3_s6_cmd_last;     
reg             m3_s6_data;         
reg             m3_s6_req_pend_tmp; 
reg             m3_s7_cmd_cur;      
reg             m3_s7_cmd_last;     
reg             m3_s7_data;         
reg             m3_s7_req_pend_tmp; 
reg             m3_s8_cmd_cur;      
reg             m3_s8_cmd_last;     
reg             m3_s8_data;         
reg             m3_s8_req_pend_tmp; 
reg             m3_s9_cmd_cur;      
reg             m3_s9_cmd_last;     
reg             m3_s9_data;         
reg             m3_s9_req_pend_tmp; 
reg     [48:0]  m4_cur_st;          
reg             m4_latch_cmd;       
reg             m4_nor_hready;      
reg     [48:0]  m4_nxt_st;          
reg             m4_s0_cmd_cur;      
reg             m4_s0_cmd_last;     
reg             m4_s0_data;         
reg             m4_s0_req_pend_tmp; 
reg             m4_s10_cmd_cur;     
reg             m4_s10_cmd_last;    
reg             m4_s10_data;        
reg             m4_s10_req_pend_tmp; 
reg             m4_s11_cmd_cur;     
reg             m4_s11_cmd_last;    
reg             m4_s11_data;        
reg             m4_s11_req_pend_tmp; 
reg             m4_s1_cmd_cur;      
reg             m4_s1_cmd_last;     
reg             m4_s1_data;         
reg             m4_s1_req_pend_tmp; 
reg             m4_s2_cmd_cur;      
reg             m4_s2_cmd_last;     
reg             m4_s2_data;         
reg             m4_s2_req_pend_tmp; 
reg             m4_s3_cmd_cur;      
reg             m4_s3_cmd_last;     
reg             m4_s3_data;         
reg             m4_s3_req_pend_tmp; 
reg             m4_s4_cmd_cur;      
reg             m4_s4_cmd_last;     
reg             m4_s4_data;         
reg             m4_s4_req_pend_tmp; 
reg             m4_s5_cmd_cur;      
reg             m4_s5_cmd_last;     
reg             m4_s5_data;         
reg             m4_s5_req_pend_tmp; 
reg             m4_s6_cmd_cur;      
reg             m4_s6_cmd_last;     
reg             m4_s6_data;         
reg             m4_s6_req_pend_tmp; 
reg             m4_s7_cmd_cur;      
reg             m4_s7_cmd_last;     
reg             m4_s7_data;         
reg             m4_s7_req_pend_tmp; 
reg             m4_s8_cmd_cur;      
reg             m4_s8_cmd_last;     
reg             m4_s8_data;         
reg             m4_s8_req_pend_tmp; 
reg             m4_s9_cmd_cur;      
reg             m4_s9_cmd_last;     
reg             m4_s9_data;         
reg             m4_s9_req_pend_tmp; 
reg     [48:0]  m5_cur_st;          
reg             m5_latch_cmd;       
reg             m5_nor_hready;      
reg     [48:0]  m5_nxt_st;          
reg             m5_s0_cmd_cur;      
reg             m5_s0_cmd_last;     
reg             m5_s0_data;         
reg             m5_s0_req_pend_tmp; 
reg             m5_s10_cmd_cur;     
reg             m5_s10_cmd_last;    
reg             m5_s10_data;        
reg             m5_s10_req_pend_tmp; 
reg             m5_s11_cmd_cur;     
reg             m5_s11_cmd_last;    
reg             m5_s11_data;        
reg             m5_s11_req_pend_tmp; 
reg             m5_s1_cmd_cur;      
reg             m5_s1_cmd_last;     
reg             m5_s1_data;         
reg             m5_s1_req_pend_tmp; 
reg             m5_s2_cmd_cur;      
reg             m5_s2_cmd_last;     
reg             m5_s2_data;         
reg             m5_s2_req_pend_tmp; 
reg             m5_s3_cmd_cur;      
reg             m5_s3_cmd_last;     
reg             m5_s3_data;         
reg             m5_s3_req_pend_tmp; 
reg             m5_s4_cmd_cur;      
reg             m5_s4_cmd_last;     
reg             m5_s4_data;         
reg             m5_s4_req_pend_tmp; 
reg             m5_s5_cmd_cur;      
reg             m5_s5_cmd_last;     
reg             m5_s5_data;         
reg             m5_s5_req_pend_tmp; 
reg             m5_s6_cmd_cur;      
reg             m5_s6_cmd_last;     
reg             m5_s6_data;         
reg             m5_s6_req_pend_tmp; 
reg             m5_s7_cmd_cur;      
reg             m5_s7_cmd_last;     
reg             m5_s7_data;         
reg             m5_s7_req_pend_tmp; 
reg             m5_s8_cmd_cur;      
reg             m5_s8_cmd_last;     
reg             m5_s8_data;         
reg             m5_s8_req_pend_tmp; 
reg             m5_s9_cmd_cur;      
reg             m5_s9_cmd_last;     
reg             m5_s9_data;         
reg             m5_s9_req_pend_tmp; 
reg     [48:0]  m6_cur_st;          
reg             m6_latch_cmd;       
reg             m6_nor_hready;      
reg     [48:0]  m6_nxt_st;          
reg             m6_s0_cmd_cur;      
reg             m6_s0_cmd_last;     
reg             m6_s0_data;         
reg             m6_s0_req_pend_tmp; 
reg             m6_s10_cmd_cur;     
reg             m6_s10_cmd_last;    
reg             m6_s10_data;        
reg             m6_s10_req_pend_tmp; 
reg             m6_s11_cmd_cur;     
reg             m6_s11_cmd_last;    
reg             m6_s11_data;        
reg             m6_s11_req_pend_tmp; 
reg             m6_s1_cmd_cur;      
reg             m6_s1_cmd_last;     
reg             m6_s1_data;         
reg             m6_s1_req_pend_tmp; 
reg             m6_s2_cmd_cur;      
reg             m6_s2_cmd_last;     
reg             m6_s2_data;         
reg             m6_s2_req_pend_tmp; 
reg             m6_s3_cmd_cur;      
reg             m6_s3_cmd_last;     
reg             m6_s3_data;         
reg             m6_s3_req_pend_tmp; 
reg             m6_s4_cmd_cur;      
reg             m6_s4_cmd_last;     
reg             m6_s4_data;         
reg             m6_s4_req_pend_tmp; 
reg             m6_s5_cmd_cur;      
reg             m6_s5_cmd_last;     
reg             m6_s5_data;         
reg             m6_s5_req_pend_tmp; 
reg             m6_s6_cmd_cur;      
reg             m6_s6_cmd_last;     
reg             m6_s6_data;         
reg             m6_s6_req_pend_tmp; 
reg             m6_s7_cmd_cur;      
reg             m6_s7_cmd_last;     
reg             m6_s7_data;         
reg             m6_s7_req_pend_tmp; 
reg             m6_s8_cmd_cur;      
reg             m6_s8_cmd_last;     
reg             m6_s8_data;         
reg             m6_s8_req_pend_tmp; 
reg             m6_s9_cmd_cur;      
reg             m6_s9_cmd_last;     
reg             m6_s9_data;         
reg             m6_s9_req_pend_tmp; 
reg     [6 :0]  s0_gnt;             
reg     [6 :0]  s10_gnt;            
reg     [6 :0]  s11_gnt;            
reg     [6 :0]  s1_gnt;             
reg     [6 :0]  s2_gnt;             
reg     [6 :0]  s3_gnt;             
reg     [6 :0]  s4_gnt;             
reg     [6 :0]  s5_gnt;             
reg     [6 :0]  s6_gnt;             
reg     [6 :0]  s7_gnt;             
reg     [6 :0]  s8_gnt;             
reg     [6 :0]  s9_gnt;             
wire            hclk;               
wire            hresetn;            
wire            m0_s0_hld;          
wire            m0_s0_req;          
wire            m0_s0_req_pend;     
wire            m0_s0_sel;          
wire            m0_s0_wt_sel;       
wire            m0_s10_hld;         
wire            m0_s10_req;         
wire            m0_s10_req_pend;    
wire            m0_s10_sel;         
wire            m0_s10_wt_sel;      
wire            m0_s11_hld;         
wire            m0_s11_req;         
wire            m0_s11_req_pend;    
wire            m0_s11_sel;         
wire            m0_s11_wt_sel;      
wire            m0_s1_hld;          
wire            m0_s1_req;          
wire            m0_s1_req_pend;     
wire            m0_s1_sel;          
wire            m0_s1_wt_sel;       
wire            m0_s2_hld;          
wire            m0_s2_req;          
wire            m0_s2_req_pend;     
wire            m0_s2_sel;          
wire            m0_s2_wt_sel;       
wire            m0_s3_hld;          
wire            m0_s3_req;          
wire            m0_s3_req_pend;     
wire            m0_s3_sel;          
wire            m0_s3_wt_sel;       
wire            m0_s4_hld;          
wire            m0_s4_req;          
wire            m0_s4_req_pend;     
wire            m0_s4_sel;          
wire            m0_s4_wt_sel;       
wire            m0_s5_hld;          
wire            m0_s5_req;          
wire            m0_s5_req_pend;     
wire            m0_s5_sel;          
wire            m0_s5_wt_sel;       
wire            m0_s6_hld;          
wire            m0_s6_req;          
wire            m0_s6_req_pend;     
wire            m0_s6_sel;          
wire            m0_s6_wt_sel;       
wire            m0_s7_hld;          
wire            m0_s7_req;          
wire            m0_s7_req_pend;     
wire            m0_s7_sel;          
wire            m0_s7_wt_sel;       
wire            m0_s8_hld;          
wire            m0_s8_req;          
wire            m0_s8_req_pend;     
wire            m0_s8_sel;          
wire            m0_s8_wt_sel;       
wire            m0_s9_hld;          
wire            m0_s9_req;          
wire            m0_s9_req_pend;     
wire            m0_s9_sel;          
wire            m0_s9_wt_sel;       
wire            m1_s0_hld;          
wire            m1_s0_req;          
wire            m1_s0_req_pend;     
wire            m1_s0_sel;          
wire            m1_s0_wt_sel;       
wire            m1_s10_hld;         
wire            m1_s10_req;         
wire            m1_s10_req_pend;    
wire            m1_s10_sel;         
wire            m1_s10_wt_sel;      
wire            m1_s11_hld;         
wire            m1_s11_req;         
wire            m1_s11_req_pend;    
wire            m1_s11_sel;         
wire            m1_s11_wt_sel;      
wire            m1_s1_hld;          
wire            m1_s1_req;          
wire            m1_s1_req_pend;     
wire            m1_s1_sel;          
wire            m1_s1_wt_sel;       
wire            m1_s2_hld;          
wire            m1_s2_req;          
wire            m1_s2_req_pend;     
wire            m1_s2_sel;          
wire            m1_s2_wt_sel;       
wire            m1_s3_hld;          
wire            m1_s3_req;          
wire            m1_s3_req_pend;     
wire            m1_s3_sel;          
wire            m1_s3_wt_sel;       
wire            m1_s4_hld;          
wire            m1_s4_req;          
wire            m1_s4_req_pend;     
wire            m1_s4_sel;          
wire            m1_s4_wt_sel;       
wire            m1_s5_hld;          
wire            m1_s5_req;          
wire            m1_s5_req_pend;     
wire            m1_s5_sel;          
wire            m1_s5_wt_sel;       
wire            m1_s6_hld;          
wire            m1_s6_req;          
wire            m1_s6_req_pend;     
wire            m1_s6_sel;          
wire            m1_s6_wt_sel;       
wire            m1_s7_hld;          
wire            m1_s7_req;          
wire            m1_s7_req_pend;     
wire            m1_s7_sel;          
wire            m1_s7_wt_sel;       
wire            m1_s8_hld;          
wire            m1_s8_req;          
wire            m1_s8_req_pend;     
wire            m1_s8_sel;          
wire            m1_s8_wt_sel;       
wire            m1_s9_hld;          
wire            m1_s9_req;          
wire            m1_s9_req_pend;     
wire            m1_s9_sel;          
wire            m1_s9_wt_sel;       
wire            m2_s0_hld;          
wire            m2_s0_req;          
wire            m2_s0_req_pend;     
wire            m2_s0_sel;          
wire            m2_s0_wt_sel;       
wire            m2_s10_hld;         
wire            m2_s10_req;         
wire            m2_s10_req_pend;    
wire            m2_s10_sel;         
wire            m2_s10_wt_sel;      
wire            m2_s11_hld;         
wire            m2_s11_req;         
wire            m2_s11_req_pend;    
wire            m2_s11_sel;         
wire            m2_s11_wt_sel;      
wire            m2_s1_hld;          
wire            m2_s1_req;          
wire            m2_s1_req_pend;     
wire            m2_s1_sel;          
wire            m2_s1_wt_sel;       
wire            m2_s2_hld;          
wire            m2_s2_req;          
wire            m2_s2_req_pend;     
wire            m2_s2_sel;          
wire            m2_s2_wt_sel;       
wire            m2_s3_hld;          
wire            m2_s3_req;          
wire            m2_s3_req_pend;     
wire            m2_s3_sel;          
wire            m2_s3_wt_sel;       
wire            m2_s4_hld;          
wire            m2_s4_req;          
wire            m2_s4_req_pend;     
wire            m2_s4_sel;          
wire            m2_s4_wt_sel;       
wire            m2_s5_hld;          
wire            m2_s5_req;          
wire            m2_s5_req_pend;     
wire            m2_s5_sel;          
wire            m2_s5_wt_sel;       
wire            m2_s6_hld;          
wire            m2_s6_req;          
wire            m2_s6_req_pend;     
wire            m2_s6_sel;          
wire            m2_s6_wt_sel;       
wire            m2_s7_hld;          
wire            m2_s7_req;          
wire            m2_s7_req_pend;     
wire            m2_s7_sel;          
wire            m2_s7_wt_sel;       
wire            m2_s8_hld;          
wire            m2_s8_req;          
wire            m2_s8_req_pend;     
wire            m2_s8_sel;          
wire            m2_s8_wt_sel;       
wire            m2_s9_hld;          
wire            m2_s9_req;          
wire            m2_s9_req_pend;     
wire            m2_s9_sel;          
wire            m2_s9_wt_sel;       
wire            m3_s0_hld;          
wire            m3_s0_req;          
wire            m3_s0_req_pend;     
wire            m3_s0_sel;          
wire            m3_s0_wt_sel;       
wire            m3_s10_hld;         
wire            m3_s10_req;         
wire            m3_s10_req_pend;    
wire            m3_s10_sel;         
wire            m3_s10_wt_sel;      
wire            m3_s11_hld;         
wire            m3_s11_req;         
wire            m3_s11_req_pend;    
wire            m3_s11_sel;         
wire            m3_s11_wt_sel;      
wire            m3_s1_hld;          
wire            m3_s1_req;          
wire            m3_s1_req_pend;     
wire            m3_s1_sel;          
wire            m3_s1_wt_sel;       
wire            m3_s2_hld;          
wire            m3_s2_req;          
wire            m3_s2_req_pend;     
wire            m3_s2_sel;          
wire            m3_s2_wt_sel;       
wire            m3_s3_hld;          
wire            m3_s3_req;          
wire            m3_s3_req_pend;     
wire            m3_s3_sel;          
wire            m3_s3_wt_sel;       
wire            m3_s4_hld;          
wire            m3_s4_req;          
wire            m3_s4_req_pend;     
wire            m3_s4_sel;          
wire            m3_s4_wt_sel;       
wire            m3_s5_hld;          
wire            m3_s5_req;          
wire            m3_s5_req_pend;     
wire            m3_s5_sel;          
wire            m3_s5_wt_sel;       
wire            m3_s6_hld;          
wire            m3_s6_req;          
wire            m3_s6_req_pend;     
wire            m3_s6_sel;          
wire            m3_s6_wt_sel;       
wire            m3_s7_hld;          
wire            m3_s7_req;          
wire            m3_s7_req_pend;     
wire            m3_s7_sel;          
wire            m3_s7_wt_sel;       
wire            m3_s8_hld;          
wire            m3_s8_req;          
wire            m3_s8_req_pend;     
wire            m3_s8_sel;          
wire            m3_s8_wt_sel;       
wire            m3_s9_hld;          
wire            m3_s9_req;          
wire            m3_s9_req_pend;     
wire            m3_s9_sel;          
wire            m3_s9_wt_sel;       
wire            m4_s0_hld;          
wire            m4_s0_req;          
wire            m4_s0_req_pend;     
wire            m4_s0_sel;          
wire            m4_s0_wt_sel;       
wire            m4_s10_hld;         
wire            m4_s10_req;         
wire            m4_s10_req_pend;    
wire            m4_s10_sel;         
wire            m4_s10_wt_sel;      
wire            m4_s11_hld;         
wire            m4_s11_req;         
wire            m4_s11_req_pend;    
wire            m4_s11_sel;         
wire            m4_s11_wt_sel;      
wire            m4_s1_hld;          
wire            m4_s1_req;          
wire            m4_s1_req_pend;     
wire            m4_s1_sel;          
wire            m4_s1_wt_sel;       
wire            m4_s2_hld;          
wire            m4_s2_req;          
wire            m4_s2_req_pend;     
wire            m4_s2_sel;          
wire            m4_s2_wt_sel;       
wire            m4_s3_hld;          
wire            m4_s3_req;          
wire            m4_s3_req_pend;     
wire            m4_s3_sel;          
wire            m4_s3_wt_sel;       
wire            m4_s4_hld;          
wire            m4_s4_req;          
wire            m4_s4_req_pend;     
wire            m4_s4_sel;          
wire            m4_s4_wt_sel;       
wire            m4_s5_hld;          
wire            m4_s5_req;          
wire            m4_s5_req_pend;     
wire            m4_s5_sel;          
wire            m4_s5_wt_sel;       
wire            m4_s6_hld;          
wire            m4_s6_req;          
wire            m4_s6_req_pend;     
wire            m4_s6_sel;          
wire            m4_s6_wt_sel;       
wire            m4_s7_hld;          
wire            m4_s7_req;          
wire            m4_s7_req_pend;     
wire            m4_s7_sel;          
wire            m4_s7_wt_sel;       
wire            m4_s8_hld;          
wire            m4_s8_req;          
wire            m4_s8_req_pend;     
wire            m4_s8_sel;          
wire            m4_s8_wt_sel;       
wire            m4_s9_hld;          
wire            m4_s9_req;          
wire            m4_s9_req_pend;     
wire            m4_s9_sel;          
wire            m4_s9_wt_sel;       
wire            m5_s0_hld;          
wire            m5_s0_req;          
wire            m5_s0_req_pend;     
wire            m5_s0_sel;          
wire            m5_s0_wt_sel;       
wire            m5_s10_hld;         
wire            m5_s10_req;         
wire            m5_s10_req_pend;    
wire            m5_s10_sel;         
wire            m5_s10_wt_sel;      
wire            m5_s11_hld;         
wire            m5_s11_req;         
wire            m5_s11_req_pend;    
wire            m5_s11_sel;         
wire            m5_s11_wt_sel;      
wire            m5_s1_hld;          
wire            m5_s1_req;          
wire            m5_s1_req_pend;     
wire            m5_s1_sel;          
wire            m5_s1_wt_sel;       
wire            m5_s2_hld;          
wire            m5_s2_req;          
wire            m5_s2_req_pend;     
wire            m5_s2_sel;          
wire            m5_s2_wt_sel;       
wire            m5_s3_hld;          
wire            m5_s3_req;          
wire            m5_s3_req_pend;     
wire            m5_s3_sel;          
wire            m5_s3_wt_sel;       
wire            m5_s4_hld;          
wire            m5_s4_req;          
wire            m5_s4_req_pend;     
wire            m5_s4_sel;          
wire            m5_s4_wt_sel;       
wire            m5_s5_hld;          
wire            m5_s5_req;          
wire            m5_s5_req_pend;     
wire            m5_s5_sel;          
wire            m5_s5_wt_sel;       
wire            m5_s6_hld;          
wire            m5_s6_req;          
wire            m5_s6_req_pend;     
wire            m5_s6_sel;          
wire            m5_s6_wt_sel;       
wire            m5_s7_hld;          
wire            m5_s7_req;          
wire            m5_s7_req_pend;     
wire            m5_s7_sel;          
wire            m5_s7_wt_sel;       
wire            m5_s8_hld;          
wire            m5_s8_req;          
wire            m5_s8_req_pend;     
wire            m5_s8_sel;          
wire            m5_s8_wt_sel;       
wire            m5_s9_hld;          
wire            m5_s9_req;          
wire            m5_s9_req_pend;     
wire            m5_s9_sel;          
wire            m5_s9_wt_sel;       
wire            m6_s0_hld;          
wire            m6_s0_req;          
wire            m6_s0_req_pend;     
wire            m6_s0_sel;          
wire            m6_s0_wt_sel;       
wire            m6_s10_hld;         
wire            m6_s10_req;         
wire            m6_s10_req_pend;    
wire            m6_s10_sel;         
wire            m6_s10_wt_sel;      
wire            m6_s11_hld;         
wire            m6_s11_req;         
wire            m6_s11_req_pend;    
wire            m6_s11_sel;         
wire            m6_s11_wt_sel;      
wire            m6_s1_hld;          
wire            m6_s1_req;          
wire            m6_s1_req_pend;     
wire            m6_s1_sel;          
wire            m6_s1_wt_sel;       
wire            m6_s2_hld;          
wire            m6_s2_req;          
wire            m6_s2_req_pend;     
wire            m6_s2_sel;          
wire            m6_s2_wt_sel;       
wire            m6_s3_hld;          
wire            m6_s3_req;          
wire            m6_s3_req_pend;     
wire            m6_s3_sel;          
wire            m6_s3_wt_sel;       
wire            m6_s4_hld;          
wire            m6_s4_req;          
wire            m6_s4_req_pend;     
wire            m6_s4_sel;          
wire            m6_s4_wt_sel;       
wire            m6_s5_hld;          
wire            m6_s5_req;          
wire            m6_s5_req_pend;     
wire            m6_s5_sel;          
wire            m6_s5_wt_sel;       
wire            m6_s6_hld;          
wire            m6_s6_req;          
wire            m6_s6_req_pend;     
wire            m6_s6_sel;          
wire            m6_s6_wt_sel;       
wire            m6_s7_hld;          
wire            m6_s7_req;          
wire            m6_s7_req_pend;     
wire            m6_s7_sel;          
wire            m6_s7_wt_sel;       
wire            m6_s8_hld;          
wire            m6_s8_req;          
wire            m6_s8_req_pend;     
wire            m6_s8_sel;          
wire            m6_s8_wt_sel;       
wire            m6_s9_hld;          
wire            m6_s9_req;          
wire            m6_s9_req_pend;     
wire            m6_s9_sel;          
wire            m6_s9_wt_sel;       
wire            s0_hready;          
wire    [6 :0]  s0_req;             
wire    [6 :0]  s0_req_all;         
wire    [6 :0]  s0_req_pend;        
wire            s10_hready;         
wire    [6 :0]  s10_req;            
wire    [6 :0]  s10_req_all;        
wire    [6 :0]  s10_req_pend;       
wire            s11_hready;         
wire    [6 :0]  s11_req;            
wire    [6 :0]  s11_req_all;        
wire    [6 :0]  s11_req_pend;       
wire            s1_hready;          
wire    [6 :0]  s1_req;             
wire    [6 :0]  s1_req_all;         
wire    [6 :0]  s1_req_pend;        
wire            s2_hready;          
wire    [6 :0]  s2_req;             
wire    [6 :0]  s2_req_all;         
wire    [6 :0]  s2_req_pend;        
wire            s3_hready;          
wire    [6 :0]  s3_req;             
wire    [6 :0]  s3_req_all;         
wire    [6 :0]  s3_req_pend;        
wire            s4_hready;          
wire    [6 :0]  s4_req;             
wire    [6 :0]  s4_req_all;         
wire    [6 :0]  s4_req_pend;        
wire            s5_hready;          
wire    [6 :0]  s5_req;             
wire    [6 :0]  s5_req_all;         
wire    [6 :0]  s5_req_pend;        
wire            s6_hready;          
wire    [6 :0]  s6_req;             
wire    [6 :0]  s6_req_all;         
wire    [6 :0]  s6_req_pend;        
wire            s7_hready;          
wire    [6 :0]  s7_req;             
wire    [6 :0]  s7_req_all;         
wire    [6 :0]  s7_req_pend;        
wire            s8_hready;          
wire    [6 :0]  s8_req;             
wire    [6 :0]  s8_req_all;         
wire    [6 :0]  s8_req_pend;        
wire            s9_hready;          
wire    [6 :0]  s9_req;             
wire    [6 :0]  s9_req_all;         
wire    [6 :0]  s9_req_pend;        
parameter S_IDLE    = 49'b0000000000000000000000000000000000000000000000001;
parameter S_S0_GNT  = 49'b0000000000000000000000000000000000000000000000010;
parameter S_S0_WAIT = 49'b0000000000000000000000000000000000000000000000100;
parameter S_S0_CMD  = 49'b0000000000000000000000000000000000000000000001000;
parameter S_S0_DATA = 49'b0000000000000000000000000000000000000000000010000;
parameter S_S1_GNT  = 49'b0000000000000000000000000000000000000000000100000;
parameter S_S1_WAIT = 49'b0000000000000000000000000000000000000000001000000;
parameter S_S1_CMD  = 49'b0000000000000000000000000000000000000000010000000;
parameter S_S1_DATA = 49'b0000000000000000000000000000000000000000100000000;
parameter S_S2_GNT  = 49'b0000000000000000000000000000000000000001000000000;
parameter S_S2_WAIT = 49'b0000000000000000000000000000000000000010000000000;
parameter S_S2_CMD  = 49'b0000000000000000000000000000000000000100000000000;
parameter S_S2_DATA = 49'b0000000000000000000000000000000000001000000000000;
parameter S_S3_GNT  = 49'b0000000000000000000000000000000000010000000000000;
parameter S_S3_WAIT = 49'b0000000000000000000000000000000000100000000000000;
parameter S_S3_CMD  = 49'b0000000000000000000000000000000001000000000000000;
parameter S_S3_DATA = 49'b0000000000000000000000000000000010000000000000000;
parameter S_S4_GNT  = 49'b0000000000000000000000000000000100000000000000000;
parameter S_S4_WAIT = 49'b0000000000000000000000000000001000000000000000000;
parameter S_S4_CMD  = 49'b0000000000000000000000000000010000000000000000000;
parameter S_S4_DATA = 49'b0000000000000000000000000000100000000000000000000;
parameter S_S5_GNT  = 49'b0000000000000000000000000001000000000000000000000;
parameter S_S5_WAIT = 49'b0000000000000000000000000010000000000000000000000;
parameter S_S5_CMD  = 49'b0000000000000000000000000100000000000000000000000;
parameter S_S5_DATA = 49'b0000000000000000000000001000000000000000000000000;
parameter S_S6_GNT  = 49'b0000000000000000000000010000000000000000000000000;
parameter S_S6_WAIT = 49'b0000000000000000000000100000000000000000000000000;
parameter S_S6_CMD  = 49'b0000000000000000000001000000000000000000000000000;
parameter S_S6_DATA = 49'b0000000000000000000010000000000000000000000000000;
parameter S_S7_GNT  = 49'b0000000000000000000100000000000000000000000000000;
parameter S_S7_WAIT = 49'b0000000000000000001000000000000000000000000000000;
parameter S_S7_CMD  = 49'b0000000000000000010000000000000000000000000000000;
parameter S_S7_DATA = 49'b0000000000000000100000000000000000000000000000000;
parameter S_S8_GNT  = 49'b0000000000000001000000000000000000000000000000000;
parameter S_S8_WAIT = 49'b0000000000000010000000000000000000000000000000000;
parameter S_S8_CMD  = 49'b0000000000000100000000000000000000000000000000000;
parameter S_S8_DATA = 49'b0000000000001000000000000000000000000000000000000;
parameter S_S9_GNT  = 49'b0000000000010000000000000000000000000000000000000;
parameter S_S9_WAIT = 49'b0000000000100000000000000000000000000000000000000;
parameter S_S9_CMD  = 49'b0000000001000000000000000000000000000000000000000;
parameter S_S9_DATA = 49'b0000000010000000000000000000000000000000000000000;
parameter S_S10_GNT  = 49'b0000000100000000000000000000000000000000000000000;
parameter S_S10_WAIT = 49'b0000001000000000000000000000000000000000000000000;
parameter S_S10_CMD  = 49'b0000010000000000000000000000000000000000000000000;
parameter S_S10_DATA = 49'b0000100000000000000000000000000000000000000000000;
parameter S_S11_GNT  = 49'b0001000000000000000000000000000000000000000000000;
parameter S_S11_WAIT = 49'b0010000000000000000000000000000000000000000000000;
parameter S_S11_CMD  = 49'b0100000000000000000000000000000000000000000000000;
parameter S_S11_DATA = 49'b1000000000000000000000000000000000000000000000000;
assign s0_req_all[7-1:0] = s0_req[7-1:0] | s0_req_pend[7-1:0];
always @( s0_req_all[6:0])
begin
casez(s0_req_all[7-1:0])
   7'b1??????: s0_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s0_gnt[7-1:0] = 7'b0100000;
   7'b001????: s0_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s0_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s0_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s0_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s0_gnt[7-1:0] = 7'b0000001;
   default: s0_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s1_req_all[7-1:0] = s1_req[7-1:0] | s1_req_pend[7-1:0];
always @( s1_req_all[6:0])
begin
casez(s1_req_all[7-1:0])
   7'b1??????: s1_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s1_gnt[7-1:0] = 7'b0100000;
   7'b001????: s1_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s1_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s1_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s1_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s1_gnt[7-1:0] = 7'b0000001;
   default: s1_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s2_req_all[7-1:0] = s2_req[7-1:0] | s2_req_pend[7-1:0];
always @( s2_req_all[6:0])
begin
casez(s2_req_all[7-1:0])
   7'b1??????: s2_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s2_gnt[7-1:0] = 7'b0100000;
   7'b001????: s2_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s2_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s2_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s2_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s2_gnt[7-1:0] = 7'b0000001;
   default: s2_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s3_req_all[7-1:0] = s3_req[7-1:0] | s3_req_pend[7-1:0];
always @( s3_req_all[6:0])
begin
casez(s3_req_all[7-1:0])
   7'b1??????: s3_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s3_gnt[7-1:0] = 7'b0100000;
   7'b001????: s3_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s3_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s3_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s3_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s3_gnt[7-1:0] = 7'b0000001;
   default: s3_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s4_req_all[7-1:0] = s4_req[7-1:0] | s4_req_pend[7-1:0];
always @( s4_req_all[6:0])
begin
casez(s4_req_all[7-1:0])
   7'b1??????: s4_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s4_gnt[7-1:0] = 7'b0100000;
   7'b001????: s4_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s4_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s4_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s4_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s4_gnt[7-1:0] = 7'b0000001;
   default: s4_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s5_req_all[7-1:0] = s5_req[7-1:0] | s5_req_pend[7-1:0];
always @( s5_req_all[6:0])
begin
casez(s5_req_all[7-1:0])
   7'b1??????: s5_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s5_gnt[7-1:0] = 7'b0100000;
   7'b001????: s5_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s5_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s5_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s5_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s5_gnt[7-1:0] = 7'b0000001;
   default: s5_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s6_req_all[7-1:0] = s6_req[7-1:0] | s6_req_pend[7-1:0];
always @( s6_req_all[6:0])
begin
casez(s6_req_all[7-1:0])
   7'b1??????: s6_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s6_gnt[7-1:0] = 7'b0100000;
   7'b001????: s6_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s6_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s6_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s6_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s6_gnt[7-1:0] = 7'b0000001;
   default: s6_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s7_req_all[7-1:0] = s7_req[7-1:0] | s7_req_pend[7-1:0];
always @( s7_req_all[6:0])
begin
casez(s7_req_all[7-1:0])
   7'b1??????: s7_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s7_gnt[7-1:0] = 7'b0100000;
   7'b001????: s7_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s7_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s7_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s7_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s7_gnt[7-1:0] = 7'b0000001;
   default: s7_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s8_req_all[7-1:0] = s8_req[7-1:0] | s8_req_pend[7-1:0];
always @( s8_req_all[6:0])
begin
casez(s8_req_all[7-1:0])
   7'b1??????: s8_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s8_gnt[7-1:0] = 7'b0100000;
   7'b001????: s8_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s8_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s8_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s8_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s8_gnt[7-1:0] = 7'b0000001;
   default: s8_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s9_req_all[7-1:0] = s9_req[7-1:0] | s9_req_pend[7-1:0];
always @( s9_req_all[6:0])
begin
casez(s9_req_all[7-1:0])
   7'b1??????: s9_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s9_gnt[7-1:0] = 7'b0100000;
   7'b001????: s9_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s9_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s9_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s9_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s9_gnt[7-1:0] = 7'b0000001;
   default: s9_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s10_req_all[7-1:0] = s10_req[7-1:0] | s10_req_pend[7-1:0];
always @( s10_req_all[6:0])
begin
casez(s10_req_all[7-1:0])
   7'b1??????: s10_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s10_gnt[7-1:0] = 7'b0100000;
   7'b001????: s10_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s10_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s10_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s10_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s10_gnt[7-1:0] = 7'b0000001;
   default: s10_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s11_req_all[7-1:0] = s11_req[7-1:0] | s11_req_pend[7-1:0];
always @( s11_req_all[6:0])
begin
casez(s11_req_all[7-1:0])
   7'b1??????: s11_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s11_gnt[7-1:0] = 7'b0100000;
   7'b001????: s11_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s11_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s11_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s11_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s11_gnt[7-1:0] = 7'b0000001;
   default: s11_gnt[7-1:0] = 7'b0000000;
endcase
end
assign m0_s0_sel = s0_gnt[6];
assign m0_s0_wt_sel = s0_req_all[6] & ~s0_gnt[6];
assign m0_s1_sel = s1_gnt[6];
assign m0_s1_wt_sel = s1_req_all[6] & ~s1_gnt[6];
assign m0_s2_sel = s2_gnt[6];
assign m0_s2_wt_sel = s2_req_all[6] & ~s2_gnt[6];
assign m0_s3_sel = s3_gnt[6];
assign m0_s3_wt_sel = s3_req_all[6] & ~s3_gnt[6];
assign m0_s4_sel = s4_gnt[6];
assign m0_s4_wt_sel = s4_req_all[6] & ~s4_gnt[6];
assign m0_s5_sel = s5_gnt[6];
assign m0_s5_wt_sel = s5_req_all[6] & ~s5_gnt[6];
assign m0_s6_sel = s6_gnt[6];
assign m0_s6_wt_sel = s6_req_all[6] & ~s6_gnt[6];
assign m0_s7_sel = s7_gnt[6];
assign m0_s7_wt_sel = s7_req_all[6] & ~s7_gnt[6];
assign m0_s8_sel = s8_gnt[6];
assign m0_s8_wt_sel = s8_req_all[6] & ~s8_gnt[6];
assign m0_s9_sel = s9_gnt[6];
assign m0_s9_wt_sel = s9_req_all[6] & ~s9_gnt[6];
assign m0_s10_sel = s10_gnt[6];
assign m0_s10_wt_sel = s10_req_all[6] & ~s10_gnt[6];
assign m0_s11_sel = s11_gnt[6];
assign m0_s11_wt_sel = s11_req_all[6] & ~s11_gnt[6];
assign m1_s0_sel = s0_gnt[5];
assign m1_s0_wt_sel = s0_req_all[5] & ~s0_gnt[5];
assign m1_s1_sel = s1_gnt[5];
assign m1_s1_wt_sel = s1_req_all[5] & ~s1_gnt[5];
assign m1_s2_sel = s2_gnt[5];
assign m1_s2_wt_sel = s2_req_all[5] & ~s2_gnt[5];
assign m1_s3_sel = s3_gnt[5];
assign m1_s3_wt_sel = s3_req_all[5] & ~s3_gnt[5];
assign m1_s4_sel = s4_gnt[5];
assign m1_s4_wt_sel = s4_req_all[5] & ~s4_gnt[5];
assign m1_s5_sel = s5_gnt[5];
assign m1_s5_wt_sel = s5_req_all[5] & ~s5_gnt[5];
assign m1_s6_sel = s6_gnt[5];
assign m1_s6_wt_sel = s6_req_all[5] & ~s6_gnt[5];
assign m1_s7_sel = s7_gnt[5];
assign m1_s7_wt_sel = s7_req_all[5] & ~s7_gnt[5];
assign m1_s8_sel = s8_gnt[5];
assign m1_s8_wt_sel = s8_req_all[5] & ~s8_gnt[5];
assign m1_s9_sel = s9_gnt[5];
assign m1_s9_wt_sel = s9_req_all[5] & ~s9_gnt[5];
assign m1_s10_sel = s10_gnt[5];
assign m1_s10_wt_sel = s10_req_all[5] & ~s10_gnt[5];
assign m1_s11_sel = s11_gnt[5];
assign m1_s11_wt_sel = s11_req_all[5] & ~s11_gnt[5];
assign m2_s0_sel = s0_gnt[4];
assign m2_s0_wt_sel = s0_req_all[4] & ~s0_gnt[4];
assign m2_s1_sel = s1_gnt[4];
assign m2_s1_wt_sel = s1_req_all[4] & ~s1_gnt[4];
assign m2_s2_sel = s2_gnt[4];
assign m2_s2_wt_sel = s2_req_all[4] & ~s2_gnt[4];
assign m2_s3_sel = s3_gnt[4];
assign m2_s3_wt_sel = s3_req_all[4] & ~s3_gnt[4];
assign m2_s4_sel = s4_gnt[4];
assign m2_s4_wt_sel = s4_req_all[4] & ~s4_gnt[4];
assign m2_s5_sel = s5_gnt[4];
assign m2_s5_wt_sel = s5_req_all[4] & ~s5_gnt[4];
assign m2_s6_sel = s6_gnt[4];
assign m2_s6_wt_sel = s6_req_all[4] & ~s6_gnt[4];
assign m2_s7_sel = s7_gnt[4];
assign m2_s7_wt_sel = s7_req_all[4] & ~s7_gnt[4];
assign m2_s8_sel = s8_gnt[4];
assign m2_s8_wt_sel = s8_req_all[4] & ~s8_gnt[4];
assign m2_s9_sel = s9_gnt[4];
assign m2_s9_wt_sel = s9_req_all[4] & ~s9_gnt[4];
assign m2_s10_sel = s10_gnt[4];
assign m2_s10_wt_sel = s10_req_all[4] & ~s10_gnt[4];
assign m2_s11_sel = s11_gnt[4];
assign m2_s11_wt_sel = s11_req_all[4] & ~s11_gnt[4];
assign m3_s0_sel = s0_gnt[3];
assign m3_s0_wt_sel = s0_req_all[3] & ~s0_gnt[3];
assign m3_s1_sel = s1_gnt[3];
assign m3_s1_wt_sel = s1_req_all[3] & ~s1_gnt[3];
assign m3_s2_sel = s2_gnt[3];
assign m3_s2_wt_sel = s2_req_all[3] & ~s2_gnt[3];
assign m3_s3_sel = s3_gnt[3];
assign m3_s3_wt_sel = s3_req_all[3] & ~s3_gnt[3];
assign m3_s4_sel = s4_gnt[3];
assign m3_s4_wt_sel = s4_req_all[3] & ~s4_gnt[3];
assign m3_s5_sel = s5_gnt[3];
assign m3_s5_wt_sel = s5_req_all[3] & ~s5_gnt[3];
assign m3_s6_sel = s6_gnt[3];
assign m3_s6_wt_sel = s6_req_all[3] & ~s6_gnt[3];
assign m3_s7_sel = s7_gnt[3];
assign m3_s7_wt_sel = s7_req_all[3] & ~s7_gnt[3];
assign m3_s8_sel = s8_gnt[3];
assign m3_s8_wt_sel = s8_req_all[3] & ~s8_gnt[3];
assign m3_s9_sel = s9_gnt[3];
assign m3_s9_wt_sel = s9_req_all[3] & ~s9_gnt[3];
assign m3_s10_sel = s10_gnt[3];
assign m3_s10_wt_sel = s10_req_all[3] & ~s10_gnt[3];
assign m3_s11_sel = s11_gnt[3];
assign m3_s11_wt_sel = s11_req_all[3] & ~s11_gnt[3];
assign m4_s0_sel = s0_gnt[2];
assign m4_s0_wt_sel = s0_req_all[2] & ~s0_gnt[2];
assign m4_s1_sel = s1_gnt[2];
assign m4_s1_wt_sel = s1_req_all[2] & ~s1_gnt[2];
assign m4_s2_sel = s2_gnt[2];
assign m4_s2_wt_sel = s2_req_all[2] & ~s2_gnt[2];
assign m4_s3_sel = s3_gnt[2];
assign m4_s3_wt_sel = s3_req_all[2] & ~s3_gnt[2];
assign m4_s4_sel = s4_gnt[2];
assign m4_s4_wt_sel = s4_req_all[2] & ~s4_gnt[2];
assign m4_s5_sel = s5_gnt[2];
assign m4_s5_wt_sel = s5_req_all[2] & ~s5_gnt[2];
assign m4_s6_sel = s6_gnt[2];
assign m4_s6_wt_sel = s6_req_all[2] & ~s6_gnt[2];
assign m4_s7_sel = s7_gnt[2];
assign m4_s7_wt_sel = s7_req_all[2] & ~s7_gnt[2];
assign m4_s8_sel = s8_gnt[2];
assign m4_s8_wt_sel = s8_req_all[2] & ~s8_gnt[2];
assign m4_s9_sel = s9_gnt[2];
assign m4_s9_wt_sel = s9_req_all[2] & ~s9_gnt[2];
assign m4_s10_sel = s10_gnt[2];
assign m4_s10_wt_sel = s10_req_all[2] & ~s10_gnt[2];
assign m4_s11_sel = s11_gnt[2];
assign m4_s11_wt_sel = s11_req_all[2] & ~s11_gnt[2];
assign m5_s0_sel = s0_gnt[1];
assign m5_s0_wt_sel = s0_req_all[1] & ~s0_gnt[1];
assign m5_s1_sel = s1_gnt[1];
assign m5_s1_wt_sel = s1_req_all[1] & ~s1_gnt[1];
assign m5_s2_sel = s2_gnt[1];
assign m5_s2_wt_sel = s2_req_all[1] & ~s2_gnt[1];
assign m5_s3_sel = s3_gnt[1];
assign m5_s3_wt_sel = s3_req_all[1] & ~s3_gnt[1];
assign m5_s4_sel = s4_gnt[1];
assign m5_s4_wt_sel = s4_req_all[1] & ~s4_gnt[1];
assign m5_s5_sel = s5_gnt[1];
assign m5_s5_wt_sel = s5_req_all[1] & ~s5_gnt[1];
assign m5_s6_sel = s6_gnt[1];
assign m5_s6_wt_sel = s6_req_all[1] & ~s6_gnt[1];
assign m5_s7_sel = s7_gnt[1];
assign m5_s7_wt_sel = s7_req_all[1] & ~s7_gnt[1];
assign m5_s8_sel = s8_gnt[1];
assign m5_s8_wt_sel = s8_req_all[1] & ~s8_gnt[1];
assign m5_s9_sel = s9_gnt[1];
assign m5_s9_wt_sel = s9_req_all[1] & ~s9_gnt[1];
assign m5_s10_sel = s10_gnt[1];
assign m5_s10_wt_sel = s10_req_all[1] & ~s10_gnt[1];
assign m5_s11_sel = s11_gnt[1];
assign m5_s11_wt_sel = s11_req_all[1] & ~s11_gnt[1];
assign m6_s0_sel = s0_gnt[0];
assign m6_s0_wt_sel = s0_req_all[0] & ~s0_gnt[0];
assign m6_s1_sel = s1_gnt[0];
assign m6_s1_wt_sel = s1_req_all[0] & ~s1_gnt[0];
assign m6_s2_sel = s2_gnt[0];
assign m6_s2_wt_sel = s2_req_all[0] & ~s2_gnt[0];
assign m6_s3_sel = s3_gnt[0];
assign m6_s3_wt_sel = s3_req_all[0] & ~s3_gnt[0];
assign m6_s4_sel = s4_gnt[0];
assign m6_s4_wt_sel = s4_req_all[0] & ~s4_gnt[0];
assign m6_s5_sel = s5_gnt[0];
assign m6_s5_wt_sel = s5_req_all[0] & ~s5_gnt[0];
assign m6_s6_sel = s6_gnt[0];
assign m6_s6_wt_sel = s6_req_all[0] & ~s6_gnt[0];
assign m6_s7_sel = s7_gnt[0];
assign m6_s7_wt_sel = s7_req_all[0] & ~s7_gnt[0];
assign m6_s8_sel = s8_gnt[0];
assign m6_s8_wt_sel = s8_req_all[0] & ~s8_gnt[0];
assign m6_s9_sel = s9_gnt[0];
assign m6_s9_wt_sel = s9_req_all[0] & ~s9_gnt[0];
assign m6_s10_sel = s10_gnt[0];
assign m6_s10_wt_sel = s10_req_all[0] & ~s10_gnt[0];
assign m6_s11_sel = s11_gnt[0];
assign m6_s11_wt_sel = s11_req_all[0] & ~s11_gnt[0];
assign m0_s0_hld =
                       (|m1_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m0_s1_hld =
                       (|m1_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m0_s2_hld =
                       (|m1_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m0_s3_hld =
                       (|m1_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m0_s4_hld =
                       (|m1_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m0_s5_hld =
                       (|m1_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m0_s6_hld =
                       (|m1_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m0_s7_hld =
                       (|m1_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m0_s8_hld =
                       (|m1_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m0_s9_hld =
                       (|m1_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m0_s10_hld =
                       (|m1_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m0_s11_hld =
                       (|m1_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m1_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m1_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m1_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m1_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m1_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m1_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m1_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m1_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m1_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m1_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m1_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m1_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m2_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m1_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m2_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m1_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m2_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m1_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m2_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m1_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m2_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m1_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m2_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m1_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m2_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m1_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m2_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m1_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m2_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m1_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m2_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m1_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m2_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m1_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m2_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m1_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m3_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m1_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m3_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m1_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m3_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m1_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m3_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m1_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m3_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m1_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m3_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m1_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m3_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m1_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m3_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m1_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m3_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m1_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m3_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m1_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m3_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m1_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m3_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m1_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m4_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m1_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m4_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m1_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m4_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m1_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m4_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m1_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m4_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m1_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m4_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m1_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m4_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m1_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m4_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m1_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m4_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m1_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m4_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m1_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m4_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m1_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m4_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m1_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m5_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m1_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m5_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m1_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m5_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m1_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m5_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m1_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m5_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m1_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m5_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m1_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m5_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m1_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m5_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m1_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m5_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m1_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m5_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m1_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m5_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m1_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m5_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m1_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m6_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m1_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]);
assign m6_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m1_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]);
assign m6_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m1_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]);
assign m6_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m1_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]);
assign m6_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m1_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]);
assign m6_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m1_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]);
assign m6_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m1_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]);
assign m6_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m1_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]);
assign m6_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m1_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]);
assign m6_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m1_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]);
assign m6_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m1_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]);
assign m6_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m1_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]);
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m0_cur_st[48:0] <= S_IDLE;
    else
       m0_cur_st[48:0] <= m0_nxt_st[48:0];
  end
always @ (*)
begin
case(m0_cur_st[48:0])
  S_IDLE:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s0_sel: begin
                          m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m0_latch_cmd = m0_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m0_s0_wt_sel: begin
                             m0_nxt_st[48:0] = S_S0_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s1_sel: begin
                          m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m0_latch_cmd = m0_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m0_s1_wt_sel: begin
                             m0_nxt_st[48:0] = S_S1_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s2_sel: begin
                          m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m0_latch_cmd = m0_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m0_s2_wt_sel: begin
                             m0_nxt_st[48:0] = S_S2_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s3_sel: begin
                          m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m0_latch_cmd = m0_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m0_s3_wt_sel: begin
                             m0_nxt_st[48:0] = S_S3_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s4_sel: begin
                          m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m0_latch_cmd = m0_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m0_s4_wt_sel: begin
                             m0_nxt_st[48:0] = S_S4_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s5_sel: begin
                          m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m0_latch_cmd = m0_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m0_s5_wt_sel: begin
                             m0_nxt_st[48:0] = S_S5_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s6_sel: begin
                          m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m0_latch_cmd = m0_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m0_s6_wt_sel: begin
                             m0_nxt_st[48:0] = S_S6_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s7_sel: begin
                          m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m0_latch_cmd = m0_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m0_s7_wt_sel: begin
                             m0_nxt_st[48:0] = S_S7_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s8_sel: begin
                          m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m0_latch_cmd = m0_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m0_s8_wt_sel: begin
                             m0_nxt_st[48:0] = S_S8_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s9_sel: begin
                          m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m0_latch_cmd = m0_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m0_s9_wt_sel: begin
                             m0_nxt_st[48:0] = S_S9_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s10_sel: begin
                          m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m0_latch_cmd = m0_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m0_s10_wt_sel: begin
                             m0_nxt_st[48:0] = S_S10_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s11_sel: begin
                          m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m0_latch_cmd = m0_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m0_s11_wt_sel: begin
                             m0_nxt_st[48:0] = S_S11_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         default: begin
                          m0_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s0_sel: begin
                          m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m0_s0_cmd_last = m0_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s1_sel: begin
                          m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m0_s1_cmd_last = m0_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s2_sel: begin
                          m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m0_s2_cmd_last = m0_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s3_sel: begin
                          m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m0_s3_cmd_last = m0_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s4_sel: begin
                          m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m0_s4_cmd_last = m0_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s5_sel: begin
                          m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m0_s5_cmd_last = m0_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s6_sel: begin
                          m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m0_s6_cmd_last = m0_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s7_sel: begin
                          m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m0_s7_cmd_last = m0_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s8_sel: begin
                          m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m0_s8_cmd_last = m0_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s9_sel: begin
                          m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m0_s9_cmd_last = m0_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s10_sel: begin
                          m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m0_s10_cmd_last = m0_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s11_sel: begin
                          m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m0_s11_cmd_last = m0_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s0_hld: begin
                          m0_nxt_st[48:0] = m0_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m0_s0_cmd_last = m0_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s1_hld: begin
                          m0_nxt_st[48:0] = m0_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m0_s1_cmd_last = m0_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s2_hld: begin
                          m0_nxt_st[48:0] = m0_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m0_s2_cmd_last = m0_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s3_hld: begin
                          m0_nxt_st[48:0] = m0_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m0_s3_cmd_last = m0_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s4_hld: begin
                          m0_nxt_st[48:0] = m0_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m0_s4_cmd_last = m0_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s5_hld: begin
                          m0_nxt_st[48:0] = m0_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m0_s5_cmd_last = m0_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s6_hld: begin
                          m0_nxt_st[48:0] = m0_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m0_s6_cmd_last = m0_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s7_hld: begin
                          m0_nxt_st[48:0] = m0_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m0_s7_cmd_last = m0_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s8_hld: begin
                          m0_nxt_st[48:0] = m0_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m0_s8_cmd_last = m0_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s9_hld: begin
                          m0_nxt_st[48:0] = m0_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m0_s9_cmd_last = m0_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s10_hld: begin
                          m0_nxt_st[48:0] = m0_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m0_s10_cmd_last = m0_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s11_hld: begin
                          m0_nxt_st[48:0] = m0_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m0_s11_cmd_last = m0_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b1;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = S_S0_DATA;
                              m0_s0_cmd_cur = 1'b1;
                             end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b1;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = S_S1_DATA;
                              m0_s1_cmd_cur = 1'b1;
                             end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b1;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = S_S2_DATA;
                              m0_s2_cmd_cur = 1'b1;
                             end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b1;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = S_S3_DATA;
                              m0_s3_cmd_cur = 1'b1;
                             end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b1;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = S_S4_DATA;
                              m0_s4_cmd_cur = 1'b1;
                             end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b1;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = S_S5_DATA;
                              m0_s5_cmd_cur = 1'b1;
                             end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b1;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = S_S6_DATA;
                              m0_s6_cmd_cur = 1'b1;
                             end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b1;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = S_S7_DATA;
                              m0_s7_cmd_cur = 1'b1;
                             end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b1;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = S_S8_DATA;
                              m0_s8_cmd_cur = 1'b1;
                             end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b1;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = S_S9_DATA;
                              m0_s9_cmd_cur = 1'b1;
                             end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b1;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = S_S10_DATA;
                              m0_s10_cmd_cur = 1'b1;
                             end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = S_S11_DATA;
                              m0_s11_cmd_cur = 1'b1;
                             end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m0_latch_cmd = 1'b0;
             m0_s0_cmd_last = 1'b0;
             m0_s0_cmd_cur = 1'b0;
             m0_s0_data = 1'b0;
             m0_s1_cmd_last = 1'b0;
             m0_s1_cmd_cur = 1'b0;
             m0_s1_data = 1'b0;
             m0_s2_cmd_last = 1'b0;
             m0_s2_cmd_cur = 1'b0;
             m0_s2_data = 1'b0;
             m0_s3_cmd_last = 1'b0;
             m0_s3_cmd_cur = 1'b0;
             m0_s3_data = 1'b0;
             m0_s4_cmd_last = 1'b0;
             m0_s4_cmd_cur = 1'b0;
             m0_s4_data = 1'b0;
             m0_s5_cmd_last = 1'b0;
             m0_s5_cmd_cur = 1'b0;
             m0_s5_data = 1'b0;
             m0_s6_cmd_last = 1'b0;
             m0_s6_cmd_cur = 1'b0;
             m0_s6_data = 1'b0;
             m0_s7_cmd_last = 1'b0;
             m0_s7_cmd_cur = 1'b0;
             m0_s7_data = 1'b0;
             m0_s8_cmd_last = 1'b0;
             m0_s8_cmd_cur = 1'b0;
             m0_s8_data = 1'b0;
             m0_s9_cmd_last = 1'b0;
             m0_s9_cmd_cur = 1'b0;
             m0_s9_data = 1'b0;
             m0_s10_cmd_last = 1'b0;
             m0_s10_cmd_cur = 1'b0;
             m0_s10_data = 1'b0;
             m0_s11_cmd_last = 1'b0;
             m0_s11_cmd_cur = 1'b0;
             m0_s11_data = 1'b0;
             m0_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m1_cur_st[48:0] <= S_IDLE;
    else
       m1_cur_st[48:0] <= m1_nxt_st[48:0];
  end
always @ (*)
begin
case(m1_cur_st[48:0])
  S_IDLE:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s0_sel: begin
                          m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m1_latch_cmd = m1_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m1_s0_wt_sel: begin
                             m1_nxt_st[48:0] = S_S0_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s1_sel: begin
                          m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m1_latch_cmd = m1_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m1_s1_wt_sel: begin
                             m1_nxt_st[48:0] = S_S1_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s2_sel: begin
                          m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m1_latch_cmd = m1_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m1_s2_wt_sel: begin
                             m1_nxt_st[48:0] = S_S2_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s3_sel: begin
                          m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m1_latch_cmd = m1_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m1_s3_wt_sel: begin
                             m1_nxt_st[48:0] = S_S3_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s4_sel: begin
                          m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m1_latch_cmd = m1_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m1_s4_wt_sel: begin
                             m1_nxt_st[48:0] = S_S4_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s5_sel: begin
                          m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m1_latch_cmd = m1_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m1_s5_wt_sel: begin
                             m1_nxt_st[48:0] = S_S5_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s6_sel: begin
                          m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m1_latch_cmd = m1_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m1_s6_wt_sel: begin
                             m1_nxt_st[48:0] = S_S6_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s7_sel: begin
                          m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m1_latch_cmd = m1_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m1_s7_wt_sel: begin
                             m1_nxt_st[48:0] = S_S7_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s8_sel: begin
                          m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m1_latch_cmd = m1_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m1_s8_wt_sel: begin
                             m1_nxt_st[48:0] = S_S8_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s9_sel: begin
                          m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m1_latch_cmd = m1_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m1_s9_wt_sel: begin
                             m1_nxt_st[48:0] = S_S9_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s10_sel: begin
                          m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m1_latch_cmd = m1_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m1_s10_wt_sel: begin
                             m1_nxt_st[48:0] = S_S10_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s11_sel: begin
                          m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m1_latch_cmd = m1_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m1_s11_wt_sel: begin
                             m1_nxt_st[48:0] = S_S11_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         default: begin
                          m1_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s0_sel: begin
                          m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m1_s0_cmd_last = m1_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s1_sel: begin
                          m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m1_s1_cmd_last = m1_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s2_sel: begin
                          m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m1_s2_cmd_last = m1_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s3_sel: begin
                          m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m1_s3_cmd_last = m1_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s4_sel: begin
                          m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m1_s4_cmd_last = m1_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s5_sel: begin
                          m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m1_s5_cmd_last = m1_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s6_sel: begin
                          m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m1_s6_cmd_last = m1_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s7_sel: begin
                          m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m1_s7_cmd_last = m1_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s8_sel: begin
                          m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m1_s8_cmd_last = m1_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s9_sel: begin
                          m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m1_s9_cmd_last = m1_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s10_sel: begin
                          m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m1_s10_cmd_last = m1_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s11_sel: begin
                          m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m1_s11_cmd_last = m1_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s0_hld: begin
                          m1_nxt_st[48:0] = m1_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m1_s0_cmd_last = m1_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s1_hld: begin
                          m1_nxt_st[48:0] = m1_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m1_s1_cmd_last = m1_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s2_hld: begin
                          m1_nxt_st[48:0] = m1_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m1_s2_cmd_last = m1_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s3_hld: begin
                          m1_nxt_st[48:0] = m1_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m1_s3_cmd_last = m1_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s4_hld: begin
                          m1_nxt_st[48:0] = m1_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m1_s4_cmd_last = m1_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s5_hld: begin
                          m1_nxt_st[48:0] = m1_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m1_s5_cmd_last = m1_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s6_hld: begin
                          m1_nxt_st[48:0] = m1_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m1_s6_cmd_last = m1_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s7_hld: begin
                          m1_nxt_st[48:0] = m1_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m1_s7_cmd_last = m1_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s8_hld: begin
                          m1_nxt_st[48:0] = m1_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m1_s8_cmd_last = m1_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s9_hld: begin
                          m1_nxt_st[48:0] = m1_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m1_s9_cmd_last = m1_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s10_hld: begin
                          m1_nxt_st[48:0] = m1_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m1_s10_cmd_last = m1_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s11_hld: begin
                          m1_nxt_st[48:0] = m1_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m1_s11_cmd_last = m1_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b1;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = S_S0_DATA;
                              m1_s0_cmd_cur = 1'b1;
                             end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b1;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = S_S1_DATA;
                              m1_s1_cmd_cur = 1'b1;
                             end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b1;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = S_S2_DATA;
                              m1_s2_cmd_cur = 1'b1;
                             end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b1;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = S_S3_DATA;
                              m1_s3_cmd_cur = 1'b1;
                             end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b1;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = S_S4_DATA;
                              m1_s4_cmd_cur = 1'b1;
                             end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b1;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = S_S5_DATA;
                              m1_s5_cmd_cur = 1'b1;
                             end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b1;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = S_S6_DATA;
                              m1_s6_cmd_cur = 1'b1;
                             end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b1;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = S_S7_DATA;
                              m1_s7_cmd_cur = 1'b1;
                             end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b1;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = S_S8_DATA;
                              m1_s8_cmd_cur = 1'b1;
                             end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b1;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = S_S9_DATA;
                              m1_s9_cmd_cur = 1'b1;
                             end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b1;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = S_S10_DATA;
                              m1_s10_cmd_cur = 1'b1;
                             end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = S_S11_DATA;
                              m1_s11_cmd_cur = 1'b1;
                             end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m1_latch_cmd = 1'b0;
             m1_s0_cmd_last = 1'b0;
             m1_s0_cmd_cur = 1'b0;
             m1_s0_data = 1'b0;
             m1_s1_cmd_last = 1'b0;
             m1_s1_cmd_cur = 1'b0;
             m1_s1_data = 1'b0;
             m1_s2_cmd_last = 1'b0;
             m1_s2_cmd_cur = 1'b0;
             m1_s2_data = 1'b0;
             m1_s3_cmd_last = 1'b0;
             m1_s3_cmd_cur = 1'b0;
             m1_s3_data = 1'b0;
             m1_s4_cmd_last = 1'b0;
             m1_s4_cmd_cur = 1'b0;
             m1_s4_data = 1'b0;
             m1_s5_cmd_last = 1'b0;
             m1_s5_cmd_cur = 1'b0;
             m1_s5_data = 1'b0;
             m1_s6_cmd_last = 1'b0;
             m1_s6_cmd_cur = 1'b0;
             m1_s6_data = 1'b0;
             m1_s7_cmd_last = 1'b0;
             m1_s7_cmd_cur = 1'b0;
             m1_s7_data = 1'b0;
             m1_s8_cmd_last = 1'b0;
             m1_s8_cmd_cur = 1'b0;
             m1_s8_data = 1'b0;
             m1_s9_cmd_last = 1'b0;
             m1_s9_cmd_cur = 1'b0;
             m1_s9_data = 1'b0;
             m1_s10_cmd_last = 1'b0;
             m1_s10_cmd_cur = 1'b0;
             m1_s10_data = 1'b0;
             m1_s11_cmd_last = 1'b0;
             m1_s11_cmd_cur = 1'b0;
             m1_s11_data = 1'b0;
             m1_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m2_cur_st[48:0] <= S_IDLE;
    else
       m2_cur_st[48:0] <= m2_nxt_st[48:0];
  end
always @ (*)
begin
case(m2_cur_st[48:0])
  S_IDLE:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s0_sel: begin
                          m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m2_latch_cmd = m2_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m2_s0_wt_sel: begin
                             m2_nxt_st[48:0] = S_S0_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s1_sel: begin
                          m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m2_latch_cmd = m2_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m2_s1_wt_sel: begin
                             m2_nxt_st[48:0] = S_S1_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s2_sel: begin
                          m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m2_latch_cmd = m2_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m2_s2_wt_sel: begin
                             m2_nxt_st[48:0] = S_S2_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s3_sel: begin
                          m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m2_latch_cmd = m2_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m2_s3_wt_sel: begin
                             m2_nxt_st[48:0] = S_S3_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s4_sel: begin
                          m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m2_latch_cmd = m2_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m2_s4_wt_sel: begin
                             m2_nxt_st[48:0] = S_S4_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s5_sel: begin
                          m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m2_latch_cmd = m2_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m2_s5_wt_sel: begin
                             m2_nxt_st[48:0] = S_S5_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s6_sel: begin
                          m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m2_latch_cmd = m2_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m2_s6_wt_sel: begin
                             m2_nxt_st[48:0] = S_S6_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s7_sel: begin
                          m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m2_latch_cmd = m2_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m2_s7_wt_sel: begin
                             m2_nxt_st[48:0] = S_S7_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s8_sel: begin
                          m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m2_latch_cmd = m2_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m2_s8_wt_sel: begin
                             m2_nxt_st[48:0] = S_S8_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s9_sel: begin
                          m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m2_latch_cmd = m2_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m2_s9_wt_sel: begin
                             m2_nxt_st[48:0] = S_S9_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s10_sel: begin
                          m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m2_latch_cmd = m2_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m2_s10_wt_sel: begin
                             m2_nxt_st[48:0] = S_S10_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s11_sel: begin
                          m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m2_latch_cmd = m2_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m2_s11_wt_sel: begin
                             m2_nxt_st[48:0] = S_S11_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         default: begin
                          m2_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s0_sel: begin
                          m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m2_s0_cmd_last = m2_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s1_sel: begin
                          m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m2_s1_cmd_last = m2_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s2_sel: begin
                          m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m2_s2_cmd_last = m2_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s3_sel: begin
                          m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m2_s3_cmd_last = m2_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s4_sel: begin
                          m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m2_s4_cmd_last = m2_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s5_sel: begin
                          m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m2_s5_cmd_last = m2_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s6_sel: begin
                          m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m2_s6_cmd_last = m2_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s7_sel: begin
                          m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m2_s7_cmd_last = m2_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s8_sel: begin
                          m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m2_s8_cmd_last = m2_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s9_sel: begin
                          m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m2_s9_cmd_last = m2_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s10_sel: begin
                          m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m2_s10_cmd_last = m2_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s11_sel: begin
                          m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m2_s11_cmd_last = m2_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s0_hld: begin
                          m2_nxt_st[48:0] = m2_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m2_s0_cmd_last = m2_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s1_hld: begin
                          m2_nxt_st[48:0] = m2_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m2_s1_cmd_last = m2_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s2_hld: begin
                          m2_nxt_st[48:0] = m2_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m2_s2_cmd_last = m2_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s3_hld: begin
                          m2_nxt_st[48:0] = m2_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m2_s3_cmd_last = m2_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s4_hld: begin
                          m2_nxt_st[48:0] = m2_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m2_s4_cmd_last = m2_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s5_hld: begin
                          m2_nxt_st[48:0] = m2_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m2_s5_cmd_last = m2_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s6_hld: begin
                          m2_nxt_st[48:0] = m2_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m2_s6_cmd_last = m2_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s7_hld: begin
                          m2_nxt_st[48:0] = m2_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m2_s7_cmd_last = m2_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s8_hld: begin
                          m2_nxt_st[48:0] = m2_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m2_s8_cmd_last = m2_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s9_hld: begin
                          m2_nxt_st[48:0] = m2_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m2_s9_cmd_last = m2_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s10_hld: begin
                          m2_nxt_st[48:0] = m2_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m2_s10_cmd_last = m2_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s11_hld: begin
                          m2_nxt_st[48:0] = m2_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m2_s11_cmd_last = m2_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b1;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = S_S0_DATA;
                              m2_s0_cmd_cur = 1'b1;
                             end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b1;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = S_S1_DATA;
                              m2_s1_cmd_cur = 1'b1;
                             end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b1;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = S_S2_DATA;
                              m2_s2_cmd_cur = 1'b1;
                             end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b1;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = S_S3_DATA;
                              m2_s3_cmd_cur = 1'b1;
                             end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b1;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = S_S4_DATA;
                              m2_s4_cmd_cur = 1'b1;
                             end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b1;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = S_S5_DATA;
                              m2_s5_cmd_cur = 1'b1;
                             end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b1;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = S_S6_DATA;
                              m2_s6_cmd_cur = 1'b1;
                             end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b1;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = S_S7_DATA;
                              m2_s7_cmd_cur = 1'b1;
                             end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b1;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = S_S8_DATA;
                              m2_s8_cmd_cur = 1'b1;
                             end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b1;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = S_S9_DATA;
                              m2_s9_cmd_cur = 1'b1;
                             end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b1;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = S_S10_DATA;
                              m2_s10_cmd_cur = 1'b1;
                             end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = S_S11_DATA;
                              m2_s11_cmd_cur = 1'b1;
                             end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m2_latch_cmd = 1'b0;
             m2_s0_cmd_last = 1'b0;
             m2_s0_cmd_cur = 1'b0;
             m2_s0_data = 1'b0;
             m2_s1_cmd_last = 1'b0;
             m2_s1_cmd_cur = 1'b0;
             m2_s1_data = 1'b0;
             m2_s2_cmd_last = 1'b0;
             m2_s2_cmd_cur = 1'b0;
             m2_s2_data = 1'b0;
             m2_s3_cmd_last = 1'b0;
             m2_s3_cmd_cur = 1'b0;
             m2_s3_data = 1'b0;
             m2_s4_cmd_last = 1'b0;
             m2_s4_cmd_cur = 1'b0;
             m2_s4_data = 1'b0;
             m2_s5_cmd_last = 1'b0;
             m2_s5_cmd_cur = 1'b0;
             m2_s5_data = 1'b0;
             m2_s6_cmd_last = 1'b0;
             m2_s6_cmd_cur = 1'b0;
             m2_s6_data = 1'b0;
             m2_s7_cmd_last = 1'b0;
             m2_s7_cmd_cur = 1'b0;
             m2_s7_data = 1'b0;
             m2_s8_cmd_last = 1'b0;
             m2_s8_cmd_cur = 1'b0;
             m2_s8_data = 1'b0;
             m2_s9_cmd_last = 1'b0;
             m2_s9_cmd_cur = 1'b0;
             m2_s9_data = 1'b0;
             m2_s10_cmd_last = 1'b0;
             m2_s10_cmd_cur = 1'b0;
             m2_s10_data = 1'b0;
             m2_s11_cmd_last = 1'b0;
             m2_s11_cmd_cur = 1'b0;
             m2_s11_data = 1'b0;
             m2_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m3_cur_st[48:0] <= S_IDLE;
    else
       m3_cur_st[48:0] <= m3_nxt_st[48:0];
  end
always @ (*)
begin
case(m3_cur_st[48:0])
  S_IDLE:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s0_sel: begin
                          m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m3_latch_cmd = m3_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m3_s0_wt_sel: begin
                             m3_nxt_st[48:0] = S_S0_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s1_sel: begin
                          m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m3_latch_cmd = m3_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m3_s1_wt_sel: begin
                             m3_nxt_st[48:0] = S_S1_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s2_sel: begin
                          m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m3_latch_cmd = m3_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m3_s2_wt_sel: begin
                             m3_nxt_st[48:0] = S_S2_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s3_sel: begin
                          m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m3_latch_cmd = m3_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m3_s3_wt_sel: begin
                             m3_nxt_st[48:0] = S_S3_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s4_sel: begin
                          m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m3_latch_cmd = m3_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m3_s4_wt_sel: begin
                             m3_nxt_st[48:0] = S_S4_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s5_sel: begin
                          m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m3_latch_cmd = m3_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m3_s5_wt_sel: begin
                             m3_nxt_st[48:0] = S_S5_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s6_sel: begin
                          m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m3_latch_cmd = m3_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m3_s6_wt_sel: begin
                             m3_nxt_st[48:0] = S_S6_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s7_sel: begin
                          m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m3_latch_cmd = m3_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m3_s7_wt_sel: begin
                             m3_nxt_st[48:0] = S_S7_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s8_sel: begin
                          m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m3_latch_cmd = m3_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m3_s8_wt_sel: begin
                             m3_nxt_st[48:0] = S_S8_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s9_sel: begin
                          m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m3_latch_cmd = m3_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m3_s9_wt_sel: begin
                             m3_nxt_st[48:0] = S_S9_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s10_sel: begin
                          m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m3_latch_cmd = m3_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m3_s10_wt_sel: begin
                             m3_nxt_st[48:0] = S_S10_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s11_sel: begin
                          m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m3_latch_cmd = m3_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m3_s11_wt_sel: begin
                             m3_nxt_st[48:0] = S_S11_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         default: begin
                          m3_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s0_sel: begin
                          m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m3_s0_cmd_last = m3_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s1_sel: begin
                          m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m3_s1_cmd_last = m3_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s2_sel: begin
                          m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m3_s2_cmd_last = m3_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s3_sel: begin
                          m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m3_s3_cmd_last = m3_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s4_sel: begin
                          m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m3_s4_cmd_last = m3_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s5_sel: begin
                          m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m3_s5_cmd_last = m3_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s6_sel: begin
                          m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m3_s6_cmd_last = m3_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s7_sel: begin
                          m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m3_s7_cmd_last = m3_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s8_sel: begin
                          m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m3_s8_cmd_last = m3_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s9_sel: begin
                          m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m3_s9_cmd_last = m3_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s10_sel: begin
                          m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m3_s10_cmd_last = m3_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s11_sel: begin
                          m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m3_s11_cmd_last = m3_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s0_hld: begin
                          m3_nxt_st[48:0] = m3_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m3_s0_cmd_last = m3_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s1_hld: begin
                          m3_nxt_st[48:0] = m3_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m3_s1_cmd_last = m3_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s2_hld: begin
                          m3_nxt_st[48:0] = m3_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m3_s2_cmd_last = m3_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s3_hld: begin
                          m3_nxt_st[48:0] = m3_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m3_s3_cmd_last = m3_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s4_hld: begin
                          m3_nxt_st[48:0] = m3_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m3_s4_cmd_last = m3_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s5_hld: begin
                          m3_nxt_st[48:0] = m3_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m3_s5_cmd_last = m3_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s6_hld: begin
                          m3_nxt_st[48:0] = m3_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m3_s6_cmd_last = m3_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s7_hld: begin
                          m3_nxt_st[48:0] = m3_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m3_s7_cmd_last = m3_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s8_hld: begin
                          m3_nxt_st[48:0] = m3_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m3_s8_cmd_last = m3_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s9_hld: begin
                          m3_nxt_st[48:0] = m3_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m3_s9_cmd_last = m3_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s10_hld: begin
                          m3_nxt_st[48:0] = m3_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m3_s10_cmd_last = m3_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s11_hld: begin
                          m3_nxt_st[48:0] = m3_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m3_s11_cmd_last = m3_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b1;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = S_S0_DATA;
                              m3_s0_cmd_cur = 1'b1;
                             end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b1;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = S_S1_DATA;
                              m3_s1_cmd_cur = 1'b1;
                             end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b1;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = S_S2_DATA;
                              m3_s2_cmd_cur = 1'b1;
                             end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b1;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = S_S3_DATA;
                              m3_s3_cmd_cur = 1'b1;
                             end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b1;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = S_S4_DATA;
                              m3_s4_cmd_cur = 1'b1;
                             end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b1;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = S_S5_DATA;
                              m3_s5_cmd_cur = 1'b1;
                             end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b1;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = S_S6_DATA;
                              m3_s6_cmd_cur = 1'b1;
                             end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b1;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = S_S7_DATA;
                              m3_s7_cmd_cur = 1'b1;
                             end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b1;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = S_S8_DATA;
                              m3_s8_cmd_cur = 1'b1;
                             end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b1;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = S_S9_DATA;
                              m3_s9_cmd_cur = 1'b1;
                             end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b1;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = S_S10_DATA;
                              m3_s10_cmd_cur = 1'b1;
                             end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = S_S11_DATA;
                              m3_s11_cmd_cur = 1'b1;
                             end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m3_latch_cmd = 1'b0;
             m3_s0_cmd_last = 1'b0;
             m3_s0_cmd_cur = 1'b0;
             m3_s0_data = 1'b0;
             m3_s1_cmd_last = 1'b0;
             m3_s1_cmd_cur = 1'b0;
             m3_s1_data = 1'b0;
             m3_s2_cmd_last = 1'b0;
             m3_s2_cmd_cur = 1'b0;
             m3_s2_data = 1'b0;
             m3_s3_cmd_last = 1'b0;
             m3_s3_cmd_cur = 1'b0;
             m3_s3_data = 1'b0;
             m3_s4_cmd_last = 1'b0;
             m3_s4_cmd_cur = 1'b0;
             m3_s4_data = 1'b0;
             m3_s5_cmd_last = 1'b0;
             m3_s5_cmd_cur = 1'b0;
             m3_s5_data = 1'b0;
             m3_s6_cmd_last = 1'b0;
             m3_s6_cmd_cur = 1'b0;
             m3_s6_data = 1'b0;
             m3_s7_cmd_last = 1'b0;
             m3_s7_cmd_cur = 1'b0;
             m3_s7_data = 1'b0;
             m3_s8_cmd_last = 1'b0;
             m3_s8_cmd_cur = 1'b0;
             m3_s8_data = 1'b0;
             m3_s9_cmd_last = 1'b0;
             m3_s9_cmd_cur = 1'b0;
             m3_s9_data = 1'b0;
             m3_s10_cmd_last = 1'b0;
             m3_s10_cmd_cur = 1'b0;
             m3_s10_data = 1'b0;
             m3_s11_cmd_last = 1'b0;
             m3_s11_cmd_cur = 1'b0;
             m3_s11_data = 1'b0;
             m3_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m4_cur_st[48:0] <= S_IDLE;
    else
       m4_cur_st[48:0] <= m4_nxt_st[48:0];
  end
always @ (*)
begin
case(m4_cur_st[48:0])
  S_IDLE:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s0_sel: begin
                          m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m4_latch_cmd = m4_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m4_s0_wt_sel: begin
                             m4_nxt_st[48:0] = S_S0_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s1_sel: begin
                          m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m4_latch_cmd = m4_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m4_s1_wt_sel: begin
                             m4_nxt_st[48:0] = S_S1_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s2_sel: begin
                          m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m4_latch_cmd = m4_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m4_s2_wt_sel: begin
                             m4_nxt_st[48:0] = S_S2_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s3_sel: begin
                          m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m4_latch_cmd = m4_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m4_s3_wt_sel: begin
                             m4_nxt_st[48:0] = S_S3_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s4_sel: begin
                          m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m4_latch_cmd = m4_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m4_s4_wt_sel: begin
                             m4_nxt_st[48:0] = S_S4_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s5_sel: begin
                          m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m4_latch_cmd = m4_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m4_s5_wt_sel: begin
                             m4_nxt_st[48:0] = S_S5_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s6_sel: begin
                          m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m4_latch_cmd = m4_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m4_s6_wt_sel: begin
                             m4_nxt_st[48:0] = S_S6_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s7_sel: begin
                          m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m4_latch_cmd = m4_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m4_s7_wt_sel: begin
                             m4_nxt_st[48:0] = S_S7_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s8_sel: begin
                          m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m4_latch_cmd = m4_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m4_s8_wt_sel: begin
                             m4_nxt_st[48:0] = S_S8_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s9_sel: begin
                          m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m4_latch_cmd = m4_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m4_s9_wt_sel: begin
                             m4_nxt_st[48:0] = S_S9_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s10_sel: begin
                          m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m4_latch_cmd = m4_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m4_s10_wt_sel: begin
                             m4_nxt_st[48:0] = S_S10_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s11_sel: begin
                          m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m4_latch_cmd = m4_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m4_s11_wt_sel: begin
                             m4_nxt_st[48:0] = S_S11_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         default: begin
                          m4_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s0_sel: begin
                          m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m4_s0_cmd_last = m4_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s1_sel: begin
                          m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m4_s1_cmd_last = m4_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s2_sel: begin
                          m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m4_s2_cmd_last = m4_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s3_sel: begin
                          m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m4_s3_cmd_last = m4_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s4_sel: begin
                          m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m4_s4_cmd_last = m4_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s5_sel: begin
                          m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m4_s5_cmd_last = m4_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s6_sel: begin
                          m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m4_s6_cmd_last = m4_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s7_sel: begin
                          m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m4_s7_cmd_last = m4_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s8_sel: begin
                          m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m4_s8_cmd_last = m4_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s9_sel: begin
                          m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m4_s9_cmd_last = m4_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s10_sel: begin
                          m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m4_s10_cmd_last = m4_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s11_sel: begin
                          m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m4_s11_cmd_last = m4_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s0_hld: begin
                          m4_nxt_st[48:0] = m4_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m4_s0_cmd_last = m4_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s1_hld: begin
                          m4_nxt_st[48:0] = m4_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m4_s1_cmd_last = m4_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s2_hld: begin
                          m4_nxt_st[48:0] = m4_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m4_s2_cmd_last = m4_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s3_hld: begin
                          m4_nxt_st[48:0] = m4_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m4_s3_cmd_last = m4_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s4_hld: begin
                          m4_nxt_st[48:0] = m4_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m4_s4_cmd_last = m4_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s5_hld: begin
                          m4_nxt_st[48:0] = m4_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m4_s5_cmd_last = m4_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s6_hld: begin
                          m4_nxt_st[48:0] = m4_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m4_s6_cmd_last = m4_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s7_hld: begin
                          m4_nxt_st[48:0] = m4_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m4_s7_cmd_last = m4_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s8_hld: begin
                          m4_nxt_st[48:0] = m4_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m4_s8_cmd_last = m4_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s9_hld: begin
                          m4_nxt_st[48:0] = m4_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m4_s9_cmd_last = m4_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s10_hld: begin
                          m4_nxt_st[48:0] = m4_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m4_s10_cmd_last = m4_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s11_hld: begin
                          m4_nxt_st[48:0] = m4_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m4_s11_cmd_last = m4_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b1;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = S_S0_DATA;
                              m4_s0_cmd_cur = 1'b1;
                             end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b1;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = S_S1_DATA;
                              m4_s1_cmd_cur = 1'b1;
                             end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b1;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = S_S2_DATA;
                              m4_s2_cmd_cur = 1'b1;
                             end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b1;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = S_S3_DATA;
                              m4_s3_cmd_cur = 1'b1;
                             end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b1;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = S_S4_DATA;
                              m4_s4_cmd_cur = 1'b1;
                             end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b1;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = S_S5_DATA;
                              m4_s5_cmd_cur = 1'b1;
                             end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b1;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = S_S6_DATA;
                              m4_s6_cmd_cur = 1'b1;
                             end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b1;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = S_S7_DATA;
                              m4_s7_cmd_cur = 1'b1;
                             end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b1;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = S_S8_DATA;
                              m4_s8_cmd_cur = 1'b1;
                             end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b1;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = S_S9_DATA;
                              m4_s9_cmd_cur = 1'b1;
                             end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b1;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = S_S10_DATA;
                              m4_s10_cmd_cur = 1'b1;
                             end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = S_S11_DATA;
                              m4_s11_cmd_cur = 1'b1;
                             end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m4_latch_cmd = 1'b0;
             m4_s0_cmd_last = 1'b0;
             m4_s0_cmd_cur = 1'b0;
             m4_s0_data = 1'b0;
             m4_s1_cmd_last = 1'b0;
             m4_s1_cmd_cur = 1'b0;
             m4_s1_data = 1'b0;
             m4_s2_cmd_last = 1'b0;
             m4_s2_cmd_cur = 1'b0;
             m4_s2_data = 1'b0;
             m4_s3_cmd_last = 1'b0;
             m4_s3_cmd_cur = 1'b0;
             m4_s3_data = 1'b0;
             m4_s4_cmd_last = 1'b0;
             m4_s4_cmd_cur = 1'b0;
             m4_s4_data = 1'b0;
             m4_s5_cmd_last = 1'b0;
             m4_s5_cmd_cur = 1'b0;
             m4_s5_data = 1'b0;
             m4_s6_cmd_last = 1'b0;
             m4_s6_cmd_cur = 1'b0;
             m4_s6_data = 1'b0;
             m4_s7_cmd_last = 1'b0;
             m4_s7_cmd_cur = 1'b0;
             m4_s7_data = 1'b0;
             m4_s8_cmd_last = 1'b0;
             m4_s8_cmd_cur = 1'b0;
             m4_s8_data = 1'b0;
             m4_s9_cmd_last = 1'b0;
             m4_s9_cmd_cur = 1'b0;
             m4_s9_data = 1'b0;
             m4_s10_cmd_last = 1'b0;
             m4_s10_cmd_cur = 1'b0;
             m4_s10_data = 1'b0;
             m4_s11_cmd_last = 1'b0;
             m4_s11_cmd_cur = 1'b0;
             m4_s11_data = 1'b0;
             m4_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m5_cur_st[48:0] <= S_IDLE;
    else
       m5_cur_st[48:0] <= m5_nxt_st[48:0];
  end
always @ (*)
begin
case(m5_cur_st[48:0])
  S_IDLE:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s0_sel: begin
                          m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m5_latch_cmd = m5_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m5_s0_wt_sel: begin
                             m5_nxt_st[48:0] = S_S0_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s1_sel: begin
                          m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m5_latch_cmd = m5_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m5_s1_wt_sel: begin
                             m5_nxt_st[48:0] = S_S1_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s2_sel: begin
                          m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m5_latch_cmd = m5_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m5_s2_wt_sel: begin
                             m5_nxt_st[48:0] = S_S2_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s3_sel: begin
                          m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m5_latch_cmd = m5_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m5_s3_wt_sel: begin
                             m5_nxt_st[48:0] = S_S3_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s4_sel: begin
                          m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m5_latch_cmd = m5_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m5_s4_wt_sel: begin
                             m5_nxt_st[48:0] = S_S4_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s5_sel: begin
                          m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m5_latch_cmd = m5_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m5_s5_wt_sel: begin
                             m5_nxt_st[48:0] = S_S5_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s6_sel: begin
                          m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m5_latch_cmd = m5_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m5_s6_wt_sel: begin
                             m5_nxt_st[48:0] = S_S6_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s7_sel: begin
                          m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m5_latch_cmd = m5_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m5_s7_wt_sel: begin
                             m5_nxt_st[48:0] = S_S7_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s8_sel: begin
                          m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m5_latch_cmd = m5_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m5_s8_wt_sel: begin
                             m5_nxt_st[48:0] = S_S8_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s9_sel: begin
                          m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m5_latch_cmd = m5_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m5_s9_wt_sel: begin
                             m5_nxt_st[48:0] = S_S9_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s10_sel: begin
                          m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m5_latch_cmd = m5_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m5_s10_wt_sel: begin
                             m5_nxt_st[48:0] = S_S10_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s11_sel: begin
                          m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m5_latch_cmd = m5_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m5_s11_wt_sel: begin
                             m5_nxt_st[48:0] = S_S11_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         default: begin
                          m5_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s0_sel: begin
                          m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m5_s0_cmd_last = m5_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s1_sel: begin
                          m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m5_s1_cmd_last = m5_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s2_sel: begin
                          m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m5_s2_cmd_last = m5_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s3_sel: begin
                          m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m5_s3_cmd_last = m5_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s4_sel: begin
                          m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m5_s4_cmd_last = m5_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s5_sel: begin
                          m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m5_s5_cmd_last = m5_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s6_sel: begin
                          m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m5_s6_cmd_last = m5_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s7_sel: begin
                          m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m5_s7_cmd_last = m5_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s8_sel: begin
                          m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m5_s8_cmd_last = m5_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s9_sel: begin
                          m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m5_s9_cmd_last = m5_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s10_sel: begin
                          m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m5_s10_cmd_last = m5_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s11_sel: begin
                          m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m5_s11_cmd_last = m5_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s0_hld: begin
                          m5_nxt_st[48:0] = m5_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m5_s0_cmd_last = m5_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s1_hld: begin
                          m5_nxt_st[48:0] = m5_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m5_s1_cmd_last = m5_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s2_hld: begin
                          m5_nxt_st[48:0] = m5_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m5_s2_cmd_last = m5_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s3_hld: begin
                          m5_nxt_st[48:0] = m5_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m5_s3_cmd_last = m5_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s4_hld: begin
                          m5_nxt_st[48:0] = m5_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m5_s4_cmd_last = m5_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s5_hld: begin
                          m5_nxt_st[48:0] = m5_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m5_s5_cmd_last = m5_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s6_hld: begin
                          m5_nxt_st[48:0] = m5_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m5_s6_cmd_last = m5_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s7_hld: begin
                          m5_nxt_st[48:0] = m5_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m5_s7_cmd_last = m5_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s8_hld: begin
                          m5_nxt_st[48:0] = m5_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m5_s8_cmd_last = m5_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s9_hld: begin
                          m5_nxt_st[48:0] = m5_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m5_s9_cmd_last = m5_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s10_hld: begin
                          m5_nxt_st[48:0] = m5_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m5_s10_cmd_last = m5_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s11_hld: begin
                          m5_nxt_st[48:0] = m5_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m5_s11_cmd_last = m5_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b1;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = S_S0_DATA;
                              m5_s0_cmd_cur = 1'b1;
                             end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b1;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = S_S1_DATA;
                              m5_s1_cmd_cur = 1'b1;
                             end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b1;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = S_S2_DATA;
                              m5_s2_cmd_cur = 1'b1;
                             end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b1;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = S_S3_DATA;
                              m5_s3_cmd_cur = 1'b1;
                             end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b1;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = S_S4_DATA;
                              m5_s4_cmd_cur = 1'b1;
                             end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b1;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = S_S5_DATA;
                              m5_s5_cmd_cur = 1'b1;
                             end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b1;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = S_S6_DATA;
                              m5_s6_cmd_cur = 1'b1;
                             end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b1;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = S_S7_DATA;
                              m5_s7_cmd_cur = 1'b1;
                             end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b1;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = S_S8_DATA;
                              m5_s8_cmd_cur = 1'b1;
                             end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b1;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = S_S9_DATA;
                              m5_s9_cmd_cur = 1'b1;
                             end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b1;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = S_S10_DATA;
                              m5_s10_cmd_cur = 1'b1;
                             end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = S_S11_DATA;
                              m5_s11_cmd_cur = 1'b1;
                             end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m5_latch_cmd = 1'b0;
             m5_s0_cmd_last = 1'b0;
             m5_s0_cmd_cur = 1'b0;
             m5_s0_data = 1'b0;
             m5_s1_cmd_last = 1'b0;
             m5_s1_cmd_cur = 1'b0;
             m5_s1_data = 1'b0;
             m5_s2_cmd_last = 1'b0;
             m5_s2_cmd_cur = 1'b0;
             m5_s2_data = 1'b0;
             m5_s3_cmd_last = 1'b0;
             m5_s3_cmd_cur = 1'b0;
             m5_s3_data = 1'b0;
             m5_s4_cmd_last = 1'b0;
             m5_s4_cmd_cur = 1'b0;
             m5_s4_data = 1'b0;
             m5_s5_cmd_last = 1'b0;
             m5_s5_cmd_cur = 1'b0;
             m5_s5_data = 1'b0;
             m5_s6_cmd_last = 1'b0;
             m5_s6_cmd_cur = 1'b0;
             m5_s6_data = 1'b0;
             m5_s7_cmd_last = 1'b0;
             m5_s7_cmd_cur = 1'b0;
             m5_s7_data = 1'b0;
             m5_s8_cmd_last = 1'b0;
             m5_s8_cmd_cur = 1'b0;
             m5_s8_data = 1'b0;
             m5_s9_cmd_last = 1'b0;
             m5_s9_cmd_cur = 1'b0;
             m5_s9_data = 1'b0;
             m5_s10_cmd_last = 1'b0;
             m5_s10_cmd_cur = 1'b0;
             m5_s10_data = 1'b0;
             m5_s11_cmd_last = 1'b0;
             m5_s11_cmd_cur = 1'b0;
             m5_s11_data = 1'b0;
             m5_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m6_cur_st[48:0] <= S_IDLE;
    else
       m6_cur_st[48:0] <= m6_nxt_st[48:0];
  end
always @ (*)
begin
case(m6_cur_st[48:0])
  S_IDLE:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s0_sel: begin
                          m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m6_latch_cmd = m6_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m6_s0_wt_sel: begin
                             m6_nxt_st[48:0] = S_S0_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s1_sel: begin
                          m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m6_latch_cmd = m6_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m6_s1_wt_sel: begin
                             m6_nxt_st[48:0] = S_S1_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s2_sel: begin
                          m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m6_latch_cmd = m6_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m6_s2_wt_sel: begin
                             m6_nxt_st[48:0] = S_S2_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s3_sel: begin
                          m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m6_latch_cmd = m6_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m6_s3_wt_sel: begin
                             m6_nxt_st[48:0] = S_S3_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s4_sel: begin
                          m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m6_latch_cmd = m6_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m6_s4_wt_sel: begin
                             m6_nxt_st[48:0] = S_S4_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s5_sel: begin
                          m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m6_latch_cmd = m6_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m6_s5_wt_sel: begin
                             m6_nxt_st[48:0] = S_S5_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s6_sel: begin
                          m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m6_latch_cmd = m6_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m6_s6_wt_sel: begin
                             m6_nxt_st[48:0] = S_S6_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s7_sel: begin
                          m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m6_latch_cmd = m6_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m6_s7_wt_sel: begin
                             m6_nxt_st[48:0] = S_S7_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s8_sel: begin
                          m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m6_latch_cmd = m6_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m6_s8_wt_sel: begin
                             m6_nxt_st[48:0] = S_S8_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s9_sel: begin
                          m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m6_latch_cmd = m6_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m6_s9_wt_sel: begin
                             m6_nxt_st[48:0] = S_S9_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s10_sel: begin
                          m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m6_latch_cmd = m6_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m6_s10_wt_sel: begin
                             m6_nxt_st[48:0] = S_S10_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s11_sel: begin
                          m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m6_latch_cmd = m6_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m6_s11_wt_sel: begin
                             m6_nxt_st[48:0] = S_S11_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         default: begin
                          m6_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s0_sel: begin
                          m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m6_s0_cmd_last = m6_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s1_sel: begin
                          m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m6_s1_cmd_last = m6_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s2_sel: begin
                          m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m6_s2_cmd_last = m6_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s3_sel: begin
                          m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m6_s3_cmd_last = m6_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s4_sel: begin
                          m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m6_s4_cmd_last = m6_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s5_sel: begin
                          m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m6_s5_cmd_last = m6_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s6_sel: begin
                          m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m6_s6_cmd_last = m6_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s7_sel: begin
                          m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m6_s7_cmd_last = m6_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s8_sel: begin
                          m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m6_s8_cmd_last = m6_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s9_sel: begin
                          m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m6_s9_cmd_last = m6_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s10_sel: begin
                          m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m6_s10_cmd_last = m6_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s11_sel: begin
                          m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m6_s11_cmd_last = m6_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s0_hld: begin
                          m6_nxt_st[48:0] = m6_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m6_s0_cmd_last = m6_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s1_hld: begin
                          m6_nxt_st[48:0] = m6_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m6_s1_cmd_last = m6_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s2_hld: begin
                          m6_nxt_st[48:0] = m6_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m6_s2_cmd_last = m6_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s3_hld: begin
                          m6_nxt_st[48:0] = m6_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m6_s3_cmd_last = m6_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s4_hld: begin
                          m6_nxt_st[48:0] = m6_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m6_s4_cmd_last = m6_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s5_hld: begin
                          m6_nxt_st[48:0] = m6_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m6_s5_cmd_last = m6_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s6_hld: begin
                          m6_nxt_st[48:0] = m6_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m6_s6_cmd_last = m6_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s7_hld: begin
                          m6_nxt_st[48:0] = m6_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m6_s7_cmd_last = m6_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s8_hld: begin
                          m6_nxt_st[48:0] = m6_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m6_s8_cmd_last = m6_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s9_hld: begin
                          m6_nxt_st[48:0] = m6_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m6_s9_cmd_last = m6_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s10_hld: begin
                          m6_nxt_st[48:0] = m6_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m6_s10_cmd_last = m6_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s11_hld: begin
                          m6_nxt_st[48:0] = m6_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m6_s11_cmd_last = m6_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b1;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = S_S0_DATA;
                              m6_s0_cmd_cur = 1'b1;
                             end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b1;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = S_S1_DATA;
                              m6_s1_cmd_cur = 1'b1;
                             end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b1;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = S_S2_DATA;
                              m6_s2_cmd_cur = 1'b1;
                             end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b1;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = S_S3_DATA;
                              m6_s3_cmd_cur = 1'b1;
                             end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b1;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = S_S4_DATA;
                              m6_s4_cmd_cur = 1'b1;
                             end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b1;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = S_S5_DATA;
                              m6_s5_cmd_cur = 1'b1;
                             end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b1;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = S_S6_DATA;
                              m6_s6_cmd_cur = 1'b1;
                             end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b1;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = S_S7_DATA;
                              m6_s7_cmd_cur = 1'b1;
                             end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b1;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = S_S8_DATA;
                              m6_s8_cmd_cur = 1'b1;
                             end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b1;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = S_S9_DATA;
                              m6_s9_cmd_cur = 1'b1;
                             end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b1;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = S_S10_DATA;
                              m6_s10_cmd_cur = 1'b1;
                             end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = S_S11_DATA;
                              m6_s11_cmd_cur = 1'b1;
                             end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m6_latch_cmd = 1'b0;
             m6_s0_cmd_last = 1'b0;
             m6_s0_cmd_cur = 1'b0;
             m6_s0_data = 1'b0;
             m6_s1_cmd_last = 1'b0;
             m6_s1_cmd_cur = 1'b0;
             m6_s1_data = 1'b0;
             m6_s2_cmd_last = 1'b0;
             m6_s2_cmd_cur = 1'b0;
             m6_s2_data = 1'b0;
             m6_s3_cmd_last = 1'b0;
             m6_s3_cmd_cur = 1'b0;
             m6_s3_data = 1'b0;
             m6_s4_cmd_last = 1'b0;
             m6_s4_cmd_cur = 1'b0;
             m6_s4_data = 1'b0;
             m6_s5_cmd_last = 1'b0;
             m6_s5_cmd_cur = 1'b0;
             m6_s5_data = 1'b0;
             m6_s6_cmd_last = 1'b0;
             m6_s6_cmd_cur = 1'b0;
             m6_s6_data = 1'b0;
             m6_s7_cmd_last = 1'b0;
             m6_s7_cmd_cur = 1'b0;
             m6_s7_data = 1'b0;
             m6_s8_cmd_last = 1'b0;
             m6_s8_cmd_cur = 1'b0;
             m6_s8_data = 1'b0;
             m6_s9_cmd_last = 1'b0;
             m6_s9_cmd_cur = 1'b0;
             m6_s9_data = 1'b0;
             m6_s10_cmd_last = 1'b0;
             m6_s10_cmd_cur = 1'b0;
             m6_s10_data = 1'b0;
             m6_s11_cmd_last = 1'b0;
             m6_s11_cmd_cur = 1'b0;
             m6_s11_data = 1'b0;
             m6_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s0_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s0_req)
        m0_s0_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m0_s0_req_pend_tmp <= 1'b0;
  end
assign m0_s0_req_pend = m0_s0_req_pend_tmp && (~((m0_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s1_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s1_req)
        m0_s1_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m0_s1_req_pend_tmp <= 1'b0;
  end
assign m0_s1_req_pend = m0_s1_req_pend_tmp && (~((m0_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s2_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s2_req)
        m0_s2_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m0_s2_req_pend_tmp <= 1'b0;
  end
assign m0_s2_req_pend = m0_s2_req_pend_tmp && (~((m0_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s3_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s3_req)
        m0_s3_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m0_s3_req_pend_tmp <= 1'b0;
  end
assign m0_s3_req_pend = m0_s3_req_pend_tmp && (~((m0_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s4_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s4_req)
        m0_s4_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m0_s4_req_pend_tmp <= 1'b0;
  end
assign m0_s4_req_pend = m0_s4_req_pend_tmp && (~((m0_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s5_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s5_req)
        m0_s5_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m0_s5_req_pend_tmp <= 1'b0;
  end
assign m0_s5_req_pend = m0_s5_req_pend_tmp && (~((m0_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s6_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s6_req)
        m0_s6_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m0_s6_req_pend_tmp <= 1'b0;
  end
assign m0_s6_req_pend = m0_s6_req_pend_tmp && (~((m0_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s7_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s7_req)
        m0_s7_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m0_s7_req_pend_tmp <= 1'b0;
  end
assign m0_s7_req_pend = m0_s7_req_pend_tmp && (~((m0_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s8_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s8_req)
        m0_s8_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m0_s8_req_pend_tmp <= 1'b0;
  end
assign m0_s8_req_pend = m0_s8_req_pend_tmp && (~((m0_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s9_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s9_req)
        m0_s9_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m0_s9_req_pend_tmp <= 1'b0;
  end
assign m0_s9_req_pend = m0_s9_req_pend_tmp && (~((m0_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s10_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s10_req)
        m0_s10_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m0_s10_req_pend_tmp <= 1'b0;
  end
assign m0_s10_req_pend = m0_s10_req_pend_tmp && (~((m0_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s11_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s11_req)
        m0_s11_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m0_s11_req_pend_tmp <= 1'b0;
  end
assign m0_s11_req_pend = m0_s11_req_pend_tmp && (~((m0_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s0_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s0_req)
        m1_s0_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m1_s0_req_pend_tmp <= 1'b0;
  end
assign m1_s0_req_pend = m1_s0_req_pend_tmp && (~((m1_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s1_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s1_req)
        m1_s1_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m1_s1_req_pend_tmp <= 1'b0;
  end
assign m1_s1_req_pend = m1_s1_req_pend_tmp && (~((m1_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s2_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s2_req)
        m1_s2_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m1_s2_req_pend_tmp <= 1'b0;
  end
assign m1_s2_req_pend = m1_s2_req_pend_tmp && (~((m1_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s3_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s3_req)
        m1_s3_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m1_s3_req_pend_tmp <= 1'b0;
  end
assign m1_s3_req_pend = m1_s3_req_pend_tmp && (~((m1_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s4_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s4_req)
        m1_s4_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m1_s4_req_pend_tmp <= 1'b0;
  end
assign m1_s4_req_pend = m1_s4_req_pend_tmp && (~((m1_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s5_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s5_req)
        m1_s5_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m1_s5_req_pend_tmp <= 1'b0;
  end
assign m1_s5_req_pend = m1_s5_req_pend_tmp && (~((m1_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s6_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s6_req)
        m1_s6_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m1_s6_req_pend_tmp <= 1'b0;
  end
assign m1_s6_req_pend = m1_s6_req_pend_tmp && (~((m1_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s7_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s7_req)
        m1_s7_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m1_s7_req_pend_tmp <= 1'b0;
  end
assign m1_s7_req_pend = m1_s7_req_pend_tmp && (~((m1_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s8_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s8_req)
        m1_s8_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m1_s8_req_pend_tmp <= 1'b0;
  end
assign m1_s8_req_pend = m1_s8_req_pend_tmp && (~((m1_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s9_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s9_req)
        m1_s9_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m1_s9_req_pend_tmp <= 1'b0;
  end
assign m1_s9_req_pend = m1_s9_req_pend_tmp && (~((m1_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s10_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s10_req)
        m1_s10_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m1_s10_req_pend_tmp <= 1'b0;
  end
assign m1_s10_req_pend = m1_s10_req_pend_tmp && (~((m1_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s11_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s11_req)
        m1_s11_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m1_s11_req_pend_tmp <= 1'b0;
  end
assign m1_s11_req_pend = m1_s11_req_pend_tmp && (~((m1_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s0_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s0_req)
        m2_s0_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m2_s0_req_pend_tmp <= 1'b0;
  end
assign m2_s0_req_pend = m2_s0_req_pend_tmp && (~((m2_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s1_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s1_req)
        m2_s1_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m2_s1_req_pend_tmp <= 1'b0;
  end
assign m2_s1_req_pend = m2_s1_req_pend_tmp && (~((m2_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s2_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s2_req)
        m2_s2_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m2_s2_req_pend_tmp <= 1'b0;
  end
assign m2_s2_req_pend = m2_s2_req_pend_tmp && (~((m2_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s3_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s3_req)
        m2_s3_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m2_s3_req_pend_tmp <= 1'b0;
  end
assign m2_s3_req_pend = m2_s3_req_pend_tmp && (~((m2_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s4_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s4_req)
        m2_s4_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m2_s4_req_pend_tmp <= 1'b0;
  end
assign m2_s4_req_pend = m2_s4_req_pend_tmp && (~((m2_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s5_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s5_req)
        m2_s5_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m2_s5_req_pend_tmp <= 1'b0;
  end
assign m2_s5_req_pend = m2_s5_req_pend_tmp && (~((m2_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s6_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s6_req)
        m2_s6_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m2_s6_req_pend_tmp <= 1'b0;
  end
assign m2_s6_req_pend = m2_s6_req_pend_tmp && (~((m2_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s7_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s7_req)
        m2_s7_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m2_s7_req_pend_tmp <= 1'b0;
  end
assign m2_s7_req_pend = m2_s7_req_pend_tmp && (~((m2_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s8_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s8_req)
        m2_s8_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m2_s8_req_pend_tmp <= 1'b0;
  end
assign m2_s8_req_pend = m2_s8_req_pend_tmp && (~((m2_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s9_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s9_req)
        m2_s9_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m2_s9_req_pend_tmp <= 1'b0;
  end
assign m2_s9_req_pend = m2_s9_req_pend_tmp && (~((m2_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s10_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s10_req)
        m2_s10_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m2_s10_req_pend_tmp <= 1'b0;
  end
assign m2_s10_req_pend = m2_s10_req_pend_tmp && (~((m2_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s11_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s11_req)
        m2_s11_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m2_s11_req_pend_tmp <= 1'b0;
  end
assign m2_s11_req_pend = m2_s11_req_pend_tmp && (~((m2_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s0_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s0_req)
        m3_s0_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m3_s0_req_pend_tmp <= 1'b0;
  end
assign m3_s0_req_pend = m3_s0_req_pend_tmp && (~((m3_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s1_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s1_req)
        m3_s1_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m3_s1_req_pend_tmp <= 1'b0;
  end
assign m3_s1_req_pend = m3_s1_req_pend_tmp && (~((m3_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s2_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s2_req)
        m3_s2_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m3_s2_req_pend_tmp <= 1'b0;
  end
assign m3_s2_req_pend = m3_s2_req_pend_tmp && (~((m3_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s3_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s3_req)
        m3_s3_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m3_s3_req_pend_tmp <= 1'b0;
  end
assign m3_s3_req_pend = m3_s3_req_pend_tmp && (~((m3_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s4_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s4_req)
        m3_s4_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m3_s4_req_pend_tmp <= 1'b0;
  end
assign m3_s4_req_pend = m3_s4_req_pend_tmp && (~((m3_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s5_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s5_req)
        m3_s5_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m3_s5_req_pend_tmp <= 1'b0;
  end
assign m3_s5_req_pend = m3_s5_req_pend_tmp && (~((m3_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s6_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s6_req)
        m3_s6_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m3_s6_req_pend_tmp <= 1'b0;
  end
assign m3_s6_req_pend = m3_s6_req_pend_tmp && (~((m3_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s7_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s7_req)
        m3_s7_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m3_s7_req_pend_tmp <= 1'b0;
  end
assign m3_s7_req_pend = m3_s7_req_pend_tmp && (~((m3_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s8_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s8_req)
        m3_s8_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m3_s8_req_pend_tmp <= 1'b0;
  end
assign m3_s8_req_pend = m3_s8_req_pend_tmp && (~((m3_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s9_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s9_req)
        m3_s9_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m3_s9_req_pend_tmp <= 1'b0;
  end
assign m3_s9_req_pend = m3_s9_req_pend_tmp && (~((m3_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s10_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s10_req)
        m3_s10_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m3_s10_req_pend_tmp <= 1'b0;
  end
assign m3_s10_req_pend = m3_s10_req_pend_tmp && (~((m3_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s11_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s11_req)
        m3_s11_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m3_s11_req_pend_tmp <= 1'b0;
  end
assign m3_s11_req_pend = m3_s11_req_pend_tmp && (~((m3_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s0_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s0_req)
        m4_s0_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m4_s0_req_pend_tmp <= 1'b0;
  end
assign m4_s0_req_pend = m4_s0_req_pend_tmp && (~((m4_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s1_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s1_req)
        m4_s1_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m4_s1_req_pend_tmp <= 1'b0;
  end
assign m4_s1_req_pend = m4_s1_req_pend_tmp && (~((m4_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s2_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s2_req)
        m4_s2_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m4_s2_req_pend_tmp <= 1'b0;
  end
assign m4_s2_req_pend = m4_s2_req_pend_tmp && (~((m4_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s3_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s3_req)
        m4_s3_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m4_s3_req_pend_tmp <= 1'b0;
  end
assign m4_s3_req_pend = m4_s3_req_pend_tmp && (~((m4_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s4_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s4_req)
        m4_s4_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m4_s4_req_pend_tmp <= 1'b0;
  end
assign m4_s4_req_pend = m4_s4_req_pend_tmp && (~((m4_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s5_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s5_req)
        m4_s5_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m4_s5_req_pend_tmp <= 1'b0;
  end
assign m4_s5_req_pend = m4_s5_req_pend_tmp && (~((m4_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s6_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s6_req)
        m4_s6_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m4_s6_req_pend_tmp <= 1'b0;
  end
assign m4_s6_req_pend = m4_s6_req_pend_tmp && (~((m4_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s7_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s7_req)
        m4_s7_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m4_s7_req_pend_tmp <= 1'b0;
  end
assign m4_s7_req_pend = m4_s7_req_pend_tmp && (~((m4_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s8_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s8_req)
        m4_s8_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m4_s8_req_pend_tmp <= 1'b0;
  end
assign m4_s8_req_pend = m4_s8_req_pend_tmp && (~((m4_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s9_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s9_req)
        m4_s9_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m4_s9_req_pend_tmp <= 1'b0;
  end
assign m4_s9_req_pend = m4_s9_req_pend_tmp && (~((m4_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s10_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s10_req)
        m4_s10_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m4_s10_req_pend_tmp <= 1'b0;
  end
assign m4_s10_req_pend = m4_s10_req_pend_tmp && (~((m4_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s11_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s11_req)
        m4_s11_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m4_s11_req_pend_tmp <= 1'b0;
  end
assign m4_s11_req_pend = m4_s11_req_pend_tmp && (~((m4_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s0_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s0_req)
        m5_s0_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m5_s0_req_pend_tmp <= 1'b0;
  end
assign m5_s0_req_pend = m5_s0_req_pend_tmp && (~((m5_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s1_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s1_req)
        m5_s1_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m5_s1_req_pend_tmp <= 1'b0;
  end
assign m5_s1_req_pend = m5_s1_req_pend_tmp && (~((m5_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s2_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s2_req)
        m5_s2_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m5_s2_req_pend_tmp <= 1'b0;
  end
assign m5_s2_req_pend = m5_s2_req_pend_tmp && (~((m5_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s3_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s3_req)
        m5_s3_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m5_s3_req_pend_tmp <= 1'b0;
  end
assign m5_s3_req_pend = m5_s3_req_pend_tmp && (~((m5_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s4_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s4_req)
        m5_s4_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m5_s4_req_pend_tmp <= 1'b0;
  end
assign m5_s4_req_pend = m5_s4_req_pend_tmp && (~((m5_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s5_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s5_req)
        m5_s5_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m5_s5_req_pend_tmp <= 1'b0;
  end
assign m5_s5_req_pend = m5_s5_req_pend_tmp && (~((m5_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s6_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s6_req)
        m5_s6_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m5_s6_req_pend_tmp <= 1'b0;
  end
assign m5_s6_req_pend = m5_s6_req_pend_tmp && (~((m5_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s7_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s7_req)
        m5_s7_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m5_s7_req_pend_tmp <= 1'b0;
  end
assign m5_s7_req_pend = m5_s7_req_pend_tmp && (~((m5_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s8_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s8_req)
        m5_s8_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m5_s8_req_pend_tmp <= 1'b0;
  end
assign m5_s8_req_pend = m5_s8_req_pend_tmp && (~((m5_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s9_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s9_req)
        m5_s9_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m5_s9_req_pend_tmp <= 1'b0;
  end
assign m5_s9_req_pend = m5_s9_req_pend_tmp && (~((m5_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s10_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s10_req)
        m5_s10_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m5_s10_req_pend_tmp <= 1'b0;
  end
assign m5_s10_req_pend = m5_s10_req_pend_tmp && (~((m5_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s11_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s11_req)
        m5_s11_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m5_s11_req_pend_tmp <= 1'b0;
  end
assign m5_s11_req_pend = m5_s11_req_pend_tmp && (~((m5_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s0_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s0_req)
        m6_s0_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m6_s0_req_pend_tmp <= 1'b0;
  end
assign m6_s0_req_pend = m6_s0_req_pend_tmp && (~((m6_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s1_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s1_req)
        m6_s1_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m6_s1_req_pend_tmp <= 1'b0;
  end
assign m6_s1_req_pend = m6_s1_req_pend_tmp && (~((m6_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s2_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s2_req)
        m6_s2_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m6_s2_req_pend_tmp <= 1'b0;
  end
assign m6_s2_req_pend = m6_s2_req_pend_tmp && (~((m6_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s3_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s3_req)
        m6_s3_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m6_s3_req_pend_tmp <= 1'b0;
  end
assign m6_s3_req_pend = m6_s3_req_pend_tmp && (~((m6_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s4_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s4_req)
        m6_s4_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m6_s4_req_pend_tmp <= 1'b0;
  end
assign m6_s4_req_pend = m6_s4_req_pend_tmp && (~((m6_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s5_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s5_req)
        m6_s5_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m6_s5_req_pend_tmp <= 1'b0;
  end
assign m6_s5_req_pend = m6_s5_req_pend_tmp && (~((m6_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s6_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s6_req)
        m6_s6_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m6_s6_req_pend_tmp <= 1'b0;
  end
assign m6_s6_req_pend = m6_s6_req_pend_tmp && (~((m6_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s7_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s7_req)
        m6_s7_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m6_s7_req_pend_tmp <= 1'b0;
  end
assign m6_s7_req_pend = m6_s7_req_pend_tmp && (~((m6_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s8_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s8_req)
        m6_s8_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m6_s8_req_pend_tmp <= 1'b0;
  end
assign m6_s8_req_pend = m6_s8_req_pend_tmp && (~((m6_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s9_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s9_req)
        m6_s9_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m6_s9_req_pend_tmp <= 1'b0;
  end
assign m6_s9_req_pend = m6_s9_req_pend_tmp && (~((m6_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s10_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s10_req)
        m6_s10_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m6_s10_req_pend_tmp <= 1'b0;
  end
assign m6_s10_req_pend = m6_s10_req_pend_tmp && (~((m6_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s11_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s11_req)
        m6_s11_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m6_s11_req_pend_tmp <= 1'b0;
  end
assign m6_s11_req_pend = m6_s11_req_pend_tmp && (~((m6_cur_st[48:0] == S_S11_DATA) && s11_hready));
assign s0_req_pend[7-1:0] = {
                        m0_s0_req_pend,
                        m1_s0_req_pend,
                        m2_s0_req_pend,
                        m3_s0_req_pend,
                        m4_s0_req_pend,
                        m5_s0_req_pend,
                        m6_s0_req_pend};
assign s1_req_pend[7-1:0] = {
                        m0_s1_req_pend,
                        m1_s1_req_pend,
                        m2_s1_req_pend,
                        m3_s1_req_pend,
                        m4_s1_req_pend,
                        m5_s1_req_pend,
                        m6_s1_req_pend};
assign s2_req_pend[7-1:0] = {
                        m0_s2_req_pend,
                        m1_s2_req_pend,
                        m2_s2_req_pend,
                        m3_s2_req_pend,
                        m4_s2_req_pend,
                        m5_s2_req_pend,
                        m6_s2_req_pend};
assign s3_req_pend[7-1:0] = {
                        m0_s3_req_pend,
                        m1_s3_req_pend,
                        m2_s3_req_pend,
                        m3_s3_req_pend,
                        m4_s3_req_pend,
                        m5_s3_req_pend,
                        m6_s3_req_pend};
assign s4_req_pend[7-1:0] = {
                        m0_s4_req_pend,
                        m1_s4_req_pend,
                        m2_s4_req_pend,
                        m3_s4_req_pend,
                        m4_s4_req_pend,
                        m5_s4_req_pend,
                        m6_s4_req_pend};
assign s5_req_pend[7-1:0] = {
                        m0_s5_req_pend,
                        m1_s5_req_pend,
                        m2_s5_req_pend,
                        m3_s5_req_pend,
                        m4_s5_req_pend,
                        m5_s5_req_pend,
                        m6_s5_req_pend};
assign s6_req_pend[7-1:0] = {
                        m0_s6_req_pend,
                        m1_s6_req_pend,
                        m2_s6_req_pend,
                        m3_s6_req_pend,
                        m4_s6_req_pend,
                        m5_s6_req_pend,
                        m6_s6_req_pend};
assign s7_req_pend[7-1:0] = {
                        m0_s7_req_pend,
                        m1_s7_req_pend,
                        m2_s7_req_pend,
                        m3_s7_req_pend,
                        m4_s7_req_pend,
                        m5_s7_req_pend,
                        m6_s7_req_pend};
assign s8_req_pend[7-1:0] = {
                        m0_s8_req_pend,
                        m1_s8_req_pend,
                        m2_s8_req_pend,
                        m3_s8_req_pend,
                        m4_s8_req_pend,
                        m5_s8_req_pend,
                        m6_s8_req_pend};
assign s9_req_pend[7-1:0] = {
                        m0_s9_req_pend,
                        m1_s9_req_pend,
                        m2_s9_req_pend,
                        m3_s9_req_pend,
                        m4_s9_req_pend,
                        m5_s9_req_pend,
                        m6_s9_req_pend};
assign s10_req_pend[7-1:0] = {
                        m0_s10_req_pend,
                        m1_s10_req_pend,
                        m2_s10_req_pend,
                        m3_s10_req_pend,
                        m4_s10_req_pend,
                        m5_s10_req_pend,
                        m6_s10_req_pend};
assign s11_req_pend[7-1:0] = {
                        m0_s11_req_pend,
                        m1_s11_req_pend,
                        m2_s11_req_pend,
                        m3_s11_req_pend,
                        m4_s11_req_pend,
                        m5_s11_req_pend,
                        m6_s11_req_pend};
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or s0_hready
       or s8_hready
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready
       or m0_cur_st[48:0])
begin
case(m0_cur_st[48:0])
   S_IDLE : m0_nor_hready = 1'b1;
   S_S0_CMD: m0_nor_hready = 1'b0;
   S_S0_GNT: m0_nor_hready = 1'b0;
   S_S0_WAIT : m0_nor_hready = 1'b0;
   S_S1_CMD: m0_nor_hready = 1'b0;
   S_S1_GNT: m0_nor_hready = 1'b0;
   S_S1_WAIT : m0_nor_hready = 1'b0;
   S_S2_CMD: m0_nor_hready = 1'b0;
   S_S2_GNT: m0_nor_hready = 1'b0;
   S_S2_WAIT : m0_nor_hready = 1'b0;
   S_S3_CMD: m0_nor_hready = 1'b0;
   S_S3_GNT: m0_nor_hready = 1'b0;
   S_S3_WAIT : m0_nor_hready = 1'b0;
   S_S4_CMD: m0_nor_hready = 1'b0;
   S_S4_GNT: m0_nor_hready = 1'b0;
   S_S4_WAIT : m0_nor_hready = 1'b0;
   S_S5_CMD: m0_nor_hready = 1'b0;
   S_S5_GNT: m0_nor_hready = 1'b0;
   S_S5_WAIT : m0_nor_hready = 1'b0;
   S_S6_CMD: m0_nor_hready = 1'b0;
   S_S6_GNT: m0_nor_hready = 1'b0;
   S_S6_WAIT : m0_nor_hready = 1'b0;
   S_S7_CMD: m0_nor_hready = 1'b0;
   S_S7_GNT: m0_nor_hready = 1'b0;
   S_S7_WAIT : m0_nor_hready = 1'b0;
   S_S8_CMD: m0_nor_hready = 1'b0;
   S_S8_GNT: m0_nor_hready = 1'b0;
   S_S8_WAIT : m0_nor_hready = 1'b0;
   S_S9_CMD: m0_nor_hready = 1'b0;
   S_S9_GNT: m0_nor_hready = 1'b0;
   S_S9_WAIT : m0_nor_hready = 1'b0;
   S_S10_CMD: m0_nor_hready = 1'b0;
   S_S10_GNT: m0_nor_hready = 1'b0;
   S_S10_WAIT : m0_nor_hready = 1'b0;
   S_S11_CMD: m0_nor_hready = 1'b0;
   S_S11_GNT: m0_nor_hready = 1'b0;
   S_S11_WAIT : m0_nor_hready = 1'b0;
   S_S0_DATA: m0_nor_hready = s0_hready;
   S_S1_DATA: m0_nor_hready = s1_hready;
   S_S2_DATA: m0_nor_hready = s2_hready;
   S_S3_DATA: m0_nor_hready = s3_hready;
   S_S4_DATA: m0_nor_hready = s4_hready;
   S_S5_DATA: m0_nor_hready = s5_hready;
   S_S6_DATA: m0_nor_hready = s6_hready;
   S_S7_DATA: m0_nor_hready = s7_hready;
   S_S8_DATA: m0_nor_hready = s8_hready;
   S_S9_DATA: m0_nor_hready = s9_hready;
   S_S10_DATA: m0_nor_hready = s10_hready;
   S_S11_DATA: m0_nor_hready = s11_hready;
   default: m0_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or m1_cur_st[48:0]
       or s0_hready
       or s8_hready
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready)
begin
case(m1_cur_st[48:0])
   S_IDLE : m1_nor_hready = 1'b1;
   S_S0_CMD: m1_nor_hready = 1'b0;
   S_S0_GNT: m1_nor_hready = 1'b0;
   S_S0_WAIT : m1_nor_hready = 1'b0;
   S_S1_CMD: m1_nor_hready = 1'b0;
   S_S1_GNT: m1_nor_hready = 1'b0;
   S_S1_WAIT : m1_nor_hready = 1'b0;
   S_S2_CMD: m1_nor_hready = 1'b0;
   S_S2_GNT: m1_nor_hready = 1'b0;
   S_S2_WAIT : m1_nor_hready = 1'b0;
   S_S3_CMD: m1_nor_hready = 1'b0;
   S_S3_GNT: m1_nor_hready = 1'b0;
   S_S3_WAIT : m1_nor_hready = 1'b0;
   S_S4_CMD: m1_nor_hready = 1'b0;
   S_S4_GNT: m1_nor_hready = 1'b0;
   S_S4_WAIT : m1_nor_hready = 1'b0;
   S_S5_CMD: m1_nor_hready = 1'b0;
   S_S5_GNT: m1_nor_hready = 1'b0;
   S_S5_WAIT : m1_nor_hready = 1'b0;
   S_S6_CMD: m1_nor_hready = 1'b0;
   S_S6_GNT: m1_nor_hready = 1'b0;
   S_S6_WAIT : m1_nor_hready = 1'b0;
   S_S7_CMD: m1_nor_hready = 1'b0;
   S_S7_GNT: m1_nor_hready = 1'b0;
   S_S7_WAIT : m1_nor_hready = 1'b0;
   S_S8_CMD: m1_nor_hready = 1'b0;
   S_S8_GNT: m1_nor_hready = 1'b0;
   S_S8_WAIT : m1_nor_hready = 1'b0;
   S_S9_CMD: m1_nor_hready = 1'b0;
   S_S9_GNT: m1_nor_hready = 1'b0;
   S_S9_WAIT : m1_nor_hready = 1'b0;
   S_S10_CMD: m1_nor_hready = 1'b0;
   S_S10_GNT: m1_nor_hready = 1'b0;
   S_S10_WAIT : m1_nor_hready = 1'b0;
   S_S11_CMD: m1_nor_hready = 1'b0;
   S_S11_GNT: m1_nor_hready = 1'b0;
   S_S11_WAIT : m1_nor_hready = 1'b0;
   S_S0_DATA: m1_nor_hready = s0_hready;
   S_S1_DATA: m1_nor_hready = s1_hready;
   S_S2_DATA: m1_nor_hready = s2_hready;
   S_S3_DATA: m1_nor_hready = s3_hready;
   S_S4_DATA: m1_nor_hready = s4_hready;
   S_S5_DATA: m1_nor_hready = s5_hready;
   S_S6_DATA: m1_nor_hready = s6_hready;
   S_S7_DATA: m1_nor_hready = s7_hready;
   S_S8_DATA: m1_nor_hready = s8_hready;
   S_S9_DATA: m1_nor_hready = s9_hready;
   S_S10_DATA: m1_nor_hready = s10_hready;
   S_S11_DATA: m1_nor_hready = s11_hready;
   default: m1_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or m2_cur_st[48:0]
       or s5_hready
       or s6_hready
       or s0_hready
       or s8_hready
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready)
begin
case(m2_cur_st[48:0])
   S_IDLE : m2_nor_hready = 1'b1;
   S_S0_CMD: m2_nor_hready = 1'b0;
   S_S0_GNT: m2_nor_hready = 1'b0;
   S_S0_WAIT : m2_nor_hready = 1'b0;
   S_S1_CMD: m2_nor_hready = 1'b0;
   S_S1_GNT: m2_nor_hready = 1'b0;
   S_S1_WAIT : m2_nor_hready = 1'b0;
   S_S2_CMD: m2_nor_hready = 1'b0;
   S_S2_GNT: m2_nor_hready = 1'b0;
   S_S2_WAIT : m2_nor_hready = 1'b0;
   S_S3_CMD: m2_nor_hready = 1'b0;
   S_S3_GNT: m2_nor_hready = 1'b0;
   S_S3_WAIT : m2_nor_hready = 1'b0;
   S_S4_CMD: m2_nor_hready = 1'b0;
   S_S4_GNT: m2_nor_hready = 1'b0;
   S_S4_WAIT : m2_nor_hready = 1'b0;
   S_S5_CMD: m2_nor_hready = 1'b0;
   S_S5_GNT: m2_nor_hready = 1'b0;
   S_S5_WAIT : m2_nor_hready = 1'b0;
   S_S6_CMD: m2_nor_hready = 1'b0;
   S_S6_GNT: m2_nor_hready = 1'b0;
   S_S6_WAIT : m2_nor_hready = 1'b0;
   S_S7_CMD: m2_nor_hready = 1'b0;
   S_S7_GNT: m2_nor_hready = 1'b0;
   S_S7_WAIT : m2_nor_hready = 1'b0;
   S_S8_CMD: m2_nor_hready = 1'b0;
   S_S8_GNT: m2_nor_hready = 1'b0;
   S_S8_WAIT : m2_nor_hready = 1'b0;
   S_S9_CMD: m2_nor_hready = 1'b0;
   S_S9_GNT: m2_nor_hready = 1'b0;
   S_S9_WAIT : m2_nor_hready = 1'b0;
   S_S10_CMD: m2_nor_hready = 1'b0;
   S_S10_GNT: m2_nor_hready = 1'b0;
   S_S10_WAIT : m2_nor_hready = 1'b0;
   S_S11_CMD: m2_nor_hready = 1'b0;
   S_S11_GNT: m2_nor_hready = 1'b0;
   S_S11_WAIT : m2_nor_hready = 1'b0;
   S_S0_DATA: m2_nor_hready = s0_hready;
   S_S1_DATA: m2_nor_hready = s1_hready;
   S_S2_DATA: m2_nor_hready = s2_hready;
   S_S3_DATA: m2_nor_hready = s3_hready;
   S_S4_DATA: m2_nor_hready = s4_hready;
   S_S5_DATA: m2_nor_hready = s5_hready;
   S_S6_DATA: m2_nor_hready = s6_hready;
   S_S7_DATA: m2_nor_hready = s7_hready;
   S_S8_DATA: m2_nor_hready = s8_hready;
   S_S9_DATA: m2_nor_hready = s9_hready;
   S_S10_DATA: m2_nor_hready = s10_hready;
   S_S11_DATA: m2_nor_hready = s11_hready;
   default: m2_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or s0_hready
       or s8_hready
       or m3_cur_st[48:0]
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready)
begin
case(m3_cur_st[48:0])
   S_IDLE : m3_nor_hready = 1'b1;
   S_S0_CMD: m3_nor_hready = 1'b0;
   S_S0_GNT: m3_nor_hready = 1'b0;
   S_S0_WAIT : m3_nor_hready = 1'b0;
   S_S1_CMD: m3_nor_hready = 1'b0;
   S_S1_GNT: m3_nor_hready = 1'b0;
   S_S1_WAIT : m3_nor_hready = 1'b0;
   S_S2_CMD: m3_nor_hready = 1'b0;
   S_S2_GNT: m3_nor_hready = 1'b0;
   S_S2_WAIT : m3_nor_hready = 1'b0;
   S_S3_CMD: m3_nor_hready = 1'b0;
   S_S3_GNT: m3_nor_hready = 1'b0;
   S_S3_WAIT : m3_nor_hready = 1'b0;
   S_S4_CMD: m3_nor_hready = 1'b0;
   S_S4_GNT: m3_nor_hready = 1'b0;
   S_S4_WAIT : m3_nor_hready = 1'b0;
   S_S5_CMD: m3_nor_hready = 1'b0;
   S_S5_GNT: m3_nor_hready = 1'b0;
   S_S5_WAIT : m3_nor_hready = 1'b0;
   S_S6_CMD: m3_nor_hready = 1'b0;
   S_S6_GNT: m3_nor_hready = 1'b0;
   S_S6_WAIT : m3_nor_hready = 1'b0;
   S_S7_CMD: m3_nor_hready = 1'b0;
   S_S7_GNT: m3_nor_hready = 1'b0;
   S_S7_WAIT : m3_nor_hready = 1'b0;
   S_S8_CMD: m3_nor_hready = 1'b0;
   S_S8_GNT: m3_nor_hready = 1'b0;
   S_S8_WAIT : m3_nor_hready = 1'b0;
   S_S9_CMD: m3_nor_hready = 1'b0;
   S_S9_GNT: m3_nor_hready = 1'b0;
   S_S9_WAIT : m3_nor_hready = 1'b0;
   S_S10_CMD: m3_nor_hready = 1'b0;
   S_S10_GNT: m3_nor_hready = 1'b0;
   S_S10_WAIT : m3_nor_hready = 1'b0;
   S_S11_CMD: m3_nor_hready = 1'b0;
   S_S11_GNT: m3_nor_hready = 1'b0;
   S_S11_WAIT : m3_nor_hready = 1'b0;
   S_S0_DATA: m3_nor_hready = s0_hready;
   S_S1_DATA: m3_nor_hready = s1_hready;
   S_S2_DATA: m3_nor_hready = s2_hready;
   S_S3_DATA: m3_nor_hready = s3_hready;
   S_S4_DATA: m3_nor_hready = s4_hready;
   S_S5_DATA: m3_nor_hready = s5_hready;
   S_S6_DATA: m3_nor_hready = s6_hready;
   S_S7_DATA: m3_nor_hready = s7_hready;
   S_S8_DATA: m3_nor_hready = s8_hready;
   S_S9_DATA: m3_nor_hready = s9_hready;
   S_S10_DATA: m3_nor_hready = s10_hready;
   S_S11_DATA: m3_nor_hready = s11_hready;
   default: m3_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or s0_hready
       or s8_hready
       or s2_hready
       or s11_hready
       or m4_cur_st[48:0]
       or s3_hready
       or s9_hready)
begin
case(m4_cur_st[48:0])
   S_IDLE : m4_nor_hready = 1'b1;
   S_S0_CMD: m4_nor_hready = 1'b0;
   S_S0_GNT: m4_nor_hready = 1'b0;
   S_S0_WAIT : m4_nor_hready = 1'b0;
   S_S1_CMD: m4_nor_hready = 1'b0;
   S_S1_GNT: m4_nor_hready = 1'b0;
   S_S1_WAIT : m4_nor_hready = 1'b0;
   S_S2_CMD: m4_nor_hready = 1'b0;
   S_S2_GNT: m4_nor_hready = 1'b0;
   S_S2_WAIT : m4_nor_hready = 1'b0;
   S_S3_CMD: m4_nor_hready = 1'b0;
   S_S3_GNT: m4_nor_hready = 1'b0;
   S_S3_WAIT : m4_nor_hready = 1'b0;
   S_S4_CMD: m4_nor_hready = 1'b0;
   S_S4_GNT: m4_nor_hready = 1'b0;
   S_S4_WAIT : m4_nor_hready = 1'b0;
   S_S5_CMD: m4_nor_hready = 1'b0;
   S_S5_GNT: m4_nor_hready = 1'b0;
   S_S5_WAIT : m4_nor_hready = 1'b0;
   S_S6_CMD: m4_nor_hready = 1'b0;
   S_S6_GNT: m4_nor_hready = 1'b0;
   S_S6_WAIT : m4_nor_hready = 1'b0;
   S_S7_CMD: m4_nor_hready = 1'b0;
   S_S7_GNT: m4_nor_hready = 1'b0;
   S_S7_WAIT : m4_nor_hready = 1'b0;
   S_S8_CMD: m4_nor_hready = 1'b0;
   S_S8_GNT: m4_nor_hready = 1'b0;
   S_S8_WAIT : m4_nor_hready = 1'b0;
   S_S9_CMD: m4_nor_hready = 1'b0;
   S_S9_GNT: m4_nor_hready = 1'b0;
   S_S9_WAIT : m4_nor_hready = 1'b0;
   S_S10_CMD: m4_nor_hready = 1'b0;
   S_S10_GNT: m4_nor_hready = 1'b0;
   S_S10_WAIT : m4_nor_hready = 1'b0;
   S_S11_CMD: m4_nor_hready = 1'b0;
   S_S11_GNT: m4_nor_hready = 1'b0;
   S_S11_WAIT : m4_nor_hready = 1'b0;
   S_S0_DATA: m4_nor_hready = s0_hready;
   S_S1_DATA: m4_nor_hready = s1_hready;
   S_S2_DATA: m4_nor_hready = s2_hready;
   S_S3_DATA: m4_nor_hready = s3_hready;
   S_S4_DATA: m4_nor_hready = s4_hready;
   S_S5_DATA: m4_nor_hready = s5_hready;
   S_S6_DATA: m4_nor_hready = s6_hready;
   S_S7_DATA: m4_nor_hready = s7_hready;
   S_S8_DATA: m4_nor_hready = s8_hready;
   S_S9_DATA: m4_nor_hready = s9_hready;
   S_S10_DATA: m4_nor_hready = s10_hready;
   S_S11_DATA: m4_nor_hready = s11_hready;
   default: m4_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or s0_hready
       or s8_hready
       or m5_cur_st[48:0]
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready)
begin
case(m5_cur_st[48:0])
   S_IDLE : m5_nor_hready = 1'b1;
   S_S0_CMD: m5_nor_hready = 1'b0;
   S_S0_GNT: m5_nor_hready = 1'b0;
   S_S0_WAIT : m5_nor_hready = 1'b0;
   S_S1_CMD: m5_nor_hready = 1'b0;
   S_S1_GNT: m5_nor_hready = 1'b0;
   S_S1_WAIT : m5_nor_hready = 1'b0;
   S_S2_CMD: m5_nor_hready = 1'b0;
   S_S2_GNT: m5_nor_hready = 1'b0;
   S_S2_WAIT : m5_nor_hready = 1'b0;
   S_S3_CMD: m5_nor_hready = 1'b0;
   S_S3_GNT: m5_nor_hready = 1'b0;
   S_S3_WAIT : m5_nor_hready = 1'b0;
   S_S4_CMD: m5_nor_hready = 1'b0;
   S_S4_GNT: m5_nor_hready = 1'b0;
   S_S4_WAIT : m5_nor_hready = 1'b0;
   S_S5_CMD: m5_nor_hready = 1'b0;
   S_S5_GNT: m5_nor_hready = 1'b0;
   S_S5_WAIT : m5_nor_hready = 1'b0;
   S_S6_CMD: m5_nor_hready = 1'b0;
   S_S6_GNT: m5_nor_hready = 1'b0;
   S_S6_WAIT : m5_nor_hready = 1'b0;
   S_S7_CMD: m5_nor_hready = 1'b0;
   S_S7_GNT: m5_nor_hready = 1'b0;
   S_S7_WAIT : m5_nor_hready = 1'b0;
   S_S8_CMD: m5_nor_hready = 1'b0;
   S_S8_GNT: m5_nor_hready = 1'b0;
   S_S8_WAIT : m5_nor_hready = 1'b0;
   S_S9_CMD: m5_nor_hready = 1'b0;
   S_S9_GNT: m5_nor_hready = 1'b0;
   S_S9_WAIT : m5_nor_hready = 1'b0;
   S_S10_CMD: m5_nor_hready = 1'b0;
   S_S10_GNT: m5_nor_hready = 1'b0;
   S_S10_WAIT : m5_nor_hready = 1'b0;
   S_S11_CMD: m5_nor_hready = 1'b0;
   S_S11_GNT: m5_nor_hready = 1'b0;
   S_S11_WAIT : m5_nor_hready = 1'b0;
   S_S0_DATA: m5_nor_hready = s0_hready;
   S_S1_DATA: m5_nor_hready = s1_hready;
   S_S2_DATA: m5_nor_hready = s2_hready;
   S_S3_DATA: m5_nor_hready = s3_hready;
   S_S4_DATA: m5_nor_hready = s4_hready;
   S_S5_DATA: m5_nor_hready = s5_hready;
   S_S6_DATA: m5_nor_hready = s6_hready;
   S_S7_DATA: m5_nor_hready = s7_hready;
   S_S8_DATA: m5_nor_hready = s8_hready;
   S_S9_DATA: m5_nor_hready = s9_hready;
   S_S10_DATA: m5_nor_hready = s10_hready;
   S_S11_DATA: m5_nor_hready = s11_hready;
   default: m5_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or m6_cur_st[48:0]
       or s0_hready
       or s8_hready
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready)
begin
case(m6_cur_st[48:0])
   S_IDLE : m6_nor_hready = 1'b1;
   S_S0_CMD: m6_nor_hready = 1'b0;
   S_S0_GNT: m6_nor_hready = 1'b0;
   S_S0_WAIT : m6_nor_hready = 1'b0;
   S_S1_CMD: m6_nor_hready = 1'b0;
   S_S1_GNT: m6_nor_hready = 1'b0;
   S_S1_WAIT : m6_nor_hready = 1'b0;
   S_S2_CMD: m6_nor_hready = 1'b0;
   S_S2_GNT: m6_nor_hready = 1'b0;
   S_S2_WAIT : m6_nor_hready = 1'b0;
   S_S3_CMD: m6_nor_hready = 1'b0;
   S_S3_GNT: m6_nor_hready = 1'b0;
   S_S3_WAIT : m6_nor_hready = 1'b0;
   S_S4_CMD: m6_nor_hready = 1'b0;
   S_S4_GNT: m6_nor_hready = 1'b0;
   S_S4_WAIT : m6_nor_hready = 1'b0;
   S_S5_CMD: m6_nor_hready = 1'b0;
   S_S5_GNT: m6_nor_hready = 1'b0;
   S_S5_WAIT : m6_nor_hready = 1'b0;
   S_S6_CMD: m6_nor_hready = 1'b0;
   S_S6_GNT: m6_nor_hready = 1'b0;
   S_S6_WAIT : m6_nor_hready = 1'b0;
   S_S7_CMD: m6_nor_hready = 1'b0;
   S_S7_GNT: m6_nor_hready = 1'b0;
   S_S7_WAIT : m6_nor_hready = 1'b0;
   S_S8_CMD: m6_nor_hready = 1'b0;
   S_S8_GNT: m6_nor_hready = 1'b0;
   S_S8_WAIT : m6_nor_hready = 1'b0;
   S_S9_CMD: m6_nor_hready = 1'b0;
   S_S9_GNT: m6_nor_hready = 1'b0;
   S_S9_WAIT : m6_nor_hready = 1'b0;
   S_S10_CMD: m6_nor_hready = 1'b0;
   S_S10_GNT: m6_nor_hready = 1'b0;
   S_S10_WAIT : m6_nor_hready = 1'b0;
   S_S11_CMD: m6_nor_hready = 1'b0;
   S_S11_GNT: m6_nor_hready = 1'b0;
   S_S11_WAIT : m6_nor_hready = 1'b0;
   S_S0_DATA: m6_nor_hready = s0_hready;
   S_S1_DATA: m6_nor_hready = s1_hready;
   S_S2_DATA: m6_nor_hready = s2_hready;
   S_S3_DATA: m6_nor_hready = s3_hready;
   S_S4_DATA: m6_nor_hready = s4_hready;
   S_S5_DATA: m6_nor_hready = s5_hready;
   S_S6_DATA: m6_nor_hready = s6_hready;
   S_S7_DATA: m6_nor_hready = s7_hready;
   S_S8_DATA: m6_nor_hready = s8_hready;
   S_S9_DATA: m6_nor_hready = s9_hready;
   S_S10_DATA: m6_nor_hready = s10_hready;
   S_S11_DATA: m6_nor_hready = s11_hready;
   default: m6_nor_hready = 1'b1;
endcase
end
endmodule
